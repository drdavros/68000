-- This file was generated with hex2rom written by Daniel Wallner

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
	port(
		A	: in std_logic_vector(11 downto 0);
		D	: out std_logic_vector(15 downto 0)
	);
end rom;

architecture rtl of rom is
begin
	process (A)
	begin
		case to_integer(unsigned(A)) is
		when 000000 => D <= "0000000000000001";	-- 0x0000
		when 000001 => D <= "0100000000000000";	-- 0x0002
		when 000002 => D <= "0000000000000000";	-- 0x0004
		when 000003 => D <= "0000010000000000";	-- 0x0006
		when 000004 => D <= "----------------";	-- 0x0008
		when 000005 => D <= "----------------";	-- 0x000A
		when 000006 => D <= "----------------";	-- 0x000C
		when 000007 => D <= "----------------";	-- 0x000E
		when 000008 => D <= "----------------";	-- 0x0010
		when 000009 => D <= "----------------";	-- 0x0012
		when 000010 => D <= "----------------";	-- 0x0014
		when 000011 => D <= "----------------";	-- 0x0016
		when 000012 => D <= "----------------";	-- 0x0018
		when 000013 => D <= "----------------";	-- 0x001A
		when 000014 => D <= "----------------";	-- 0x001C
		when 000015 => D <= "----------------";	-- 0x001E
		when 000016 => D <= "----------------";	-- 0x0020
		when 000017 => D <= "----------------";	-- 0x0022
		when 000018 => D <= "----------------";	-- 0x0024
		when 000019 => D <= "----------------";	-- 0x0026
		when 000020 => D <= "----------------";	-- 0x0028
		when 000021 => D <= "----------------";	-- 0x002A
		when 000022 => D <= "----------------";	-- 0x002C
		when 000023 => D <= "----------------";	-- 0x002E
		when 000024 => D <= "----------------";	-- 0x0030
		when 000025 => D <= "----------------";	-- 0x0032
		when 000026 => D <= "----------------";	-- 0x0034
		when 000027 => D <= "----------------";	-- 0x0036
		when 000028 => D <= "----------------";	-- 0x0038
		when 000029 => D <= "----------------";	-- 0x003A
		when 000030 => D <= "----------------";	-- 0x003C
		when 000031 => D <= "----------------";	-- 0x003E
		when 000032 => D <= "----------------";	-- 0x0040
		when 000033 => D <= "----------------";	-- 0x0042
		when 000034 => D <= "----------------";	-- 0x0044
		when 000035 => D <= "----------------";	-- 0x0046
		when 000036 => D <= "----------------";	-- 0x0048
		when 000037 => D <= "----------------";	-- 0x004A
		when 000038 => D <= "----------------";	-- 0x004C
		when 000039 => D <= "----------------";	-- 0x004E
		when 000040 => D <= "----------------";	-- 0x0050
		when 000041 => D <= "----------------";	-- 0x0052
		when 000042 => D <= "----------------";	-- 0x0054
		when 000043 => D <= "----------------";	-- 0x0056
		when 000044 => D <= "----------------";	-- 0x0058
		when 000045 => D <= "----------------";	-- 0x005A
		when 000046 => D <= "----------------";	-- 0x005C
		when 000047 => D <= "----------------";	-- 0x005E
		when 000048 => D <= "----------------";	-- 0x0060
		when 000049 => D <= "----------------";	-- 0x0062
		when 000050 => D <= "----------------";	-- 0x0064
		when 000051 => D <= "----------------";	-- 0x0066
		when 000052 => D <= "----------------";	-- 0x0068
		when 000053 => D <= "----------------";	-- 0x006A
		when 000054 => D <= "----------------";	-- 0x006C
		when 000055 => D <= "----------------";	-- 0x006E
		when 000056 => D <= "----------------";	-- 0x0070
		when 000057 => D <= "----------------";	-- 0x0072
		when 000058 => D <= "----------------";	-- 0x0074
		when 000059 => D <= "----------------";	-- 0x0076
		when 000060 => D <= "----------------";	-- 0x0078
		when 000061 => D <= "----------------";	-- 0x007A
		when 000062 => D <= "----------------";	-- 0x007C
		when 000063 => D <= "----------------";	-- 0x007E
		when 000064 => D <= "----------------";	-- 0x0080
		when 000065 => D <= "----------------";	-- 0x0082
		when 000066 => D <= "----------------";	-- 0x0084
		when 000067 => D <= "----------------";	-- 0x0086
		when 000068 => D <= "----------------";	-- 0x0088
		when 000069 => D <= "----------------";	-- 0x008A
		when 000070 => D <= "----------------";	-- 0x008C
		when 000071 => D <= "----------------";	-- 0x008E
		when 000072 => D <= "----------------";	-- 0x0090
		when 000073 => D <= "----------------";	-- 0x0092
		when 000074 => D <= "----------------";	-- 0x0094
		when 000075 => D <= "----------------";	-- 0x0096
		when 000076 => D <= "----------------";	-- 0x0098
		when 000077 => D <= "----------------";	-- 0x009A
		when 000078 => D <= "----------------";	-- 0x009C
		when 000079 => D <= "----------------";	-- 0x009E
		when 000080 => D <= "----------------";	-- 0x00A0
		when 000081 => D <= "----------------";	-- 0x00A2
		when 000082 => D <= "----------------";	-- 0x00A4
		when 000083 => D <= "----------------";	-- 0x00A6
		when 000084 => D <= "----------------";	-- 0x00A8
		when 000085 => D <= "----------------";	-- 0x00AA
		when 000086 => D <= "----------------";	-- 0x00AC
		when 000087 => D <= "----------------";	-- 0x00AE
		when 000088 => D <= "----------------";	-- 0x00B0
		when 000089 => D <= "----------------";	-- 0x00B2
		when 000090 => D <= "----------------";	-- 0x00B4
		when 000091 => D <= "----------------";	-- 0x00B6
		when 000092 => D <= "----------------";	-- 0x00B8
		when 000093 => D <= "----------------";	-- 0x00BA
		when 000094 => D <= "----------------";	-- 0x00BC
		when 000095 => D <= "----------------";	-- 0x00BE
		when 000096 => D <= "----------------";	-- 0x00C0
		when 000097 => D <= "----------------";	-- 0x00C2
		when 000098 => D <= "----------------";	-- 0x00C4
		when 000099 => D <= "----------------";	-- 0x00C6
		when 000100 => D <= "----------------";	-- 0x00C8
		when 000101 => D <= "----------------";	-- 0x00CA
		when 000102 => D <= "----------------";	-- 0x00CC
		when 000103 => D <= "----------------";	-- 0x00CE
		when 000104 => D <= "----------------";	-- 0x00D0
		when 000105 => D <= "----------------";	-- 0x00D2
		when 000106 => D <= "----------------";	-- 0x00D4
		when 000107 => D <= "----------------";	-- 0x00D6
		when 000108 => D <= "----------------";	-- 0x00D8
		when 000109 => D <= "----------------";	-- 0x00DA
		when 000110 => D <= "----------------";	-- 0x00DC
		when 000111 => D <= "----------------";	-- 0x00DE
		when 000112 => D <= "----------------";	-- 0x00E0
		when 000113 => D <= "----------------";	-- 0x00E2
		when 000114 => D <= "----------------";	-- 0x00E4
		when 000115 => D <= "----------------";	-- 0x00E6
		when 000116 => D <= "----------------";	-- 0x00E8
		when 000117 => D <= "----------------";	-- 0x00EA
		when 000118 => D <= "----------------";	-- 0x00EC
		when 000119 => D <= "----------------";	-- 0x00EE
		when 000120 => D <= "----------------";	-- 0x00F0
		when 000121 => D <= "----------------";	-- 0x00F2
		when 000122 => D <= "----------------";	-- 0x00F4
		when 000123 => D <= "----------------";	-- 0x00F6
		when 000124 => D <= "----------------";	-- 0x00F8
		when 000125 => D <= "----------------";	-- 0x00FA
		when 000126 => D <= "----------------";	-- 0x00FC
		when 000127 => D <= "----------------";	-- 0x00FE
		when 000128 => D <= "----------------";	-- 0x0100
		when 000129 => D <= "----------------";	-- 0x0102
		when 000130 => D <= "----------------";	-- 0x0104
		when 000131 => D <= "----------------";	-- 0x0106
		when 000132 => D <= "----------------";	-- 0x0108
		when 000133 => D <= "----------------";	-- 0x010A
		when 000134 => D <= "----------------";	-- 0x010C
		when 000135 => D <= "----------------";	-- 0x010E
		when 000136 => D <= "----------------";	-- 0x0110
		when 000137 => D <= "----------------";	-- 0x0112
		when 000138 => D <= "----------------";	-- 0x0114
		when 000139 => D <= "----------------";	-- 0x0116
		when 000140 => D <= "----------------";	-- 0x0118
		when 000141 => D <= "----------------";	-- 0x011A
		when 000142 => D <= "----------------";	-- 0x011C
		when 000143 => D <= "----------------";	-- 0x011E
		when 000144 => D <= "----------------";	-- 0x0120
		when 000145 => D <= "----------------";	-- 0x0122
		when 000146 => D <= "----------------";	-- 0x0124
		when 000147 => D <= "----------------";	-- 0x0126
		when 000148 => D <= "----------------";	-- 0x0128
		when 000149 => D <= "----------------";	-- 0x012A
		when 000150 => D <= "----------------";	-- 0x012C
		when 000151 => D <= "----------------";	-- 0x012E
		when 000152 => D <= "----------------";	-- 0x0130
		when 000153 => D <= "----------------";	-- 0x0132
		when 000154 => D <= "----------------";	-- 0x0134
		when 000155 => D <= "----------------";	-- 0x0136
		when 000156 => D <= "----------------";	-- 0x0138
		when 000157 => D <= "----------------";	-- 0x013A
		when 000158 => D <= "----------------";	-- 0x013C
		when 000159 => D <= "----------------";	-- 0x013E
		when 000160 => D <= "----------------";	-- 0x0140
		when 000161 => D <= "----------------";	-- 0x0142
		when 000162 => D <= "----------------";	-- 0x0144
		when 000163 => D <= "----------------";	-- 0x0146
		when 000164 => D <= "----------------";	-- 0x0148
		when 000165 => D <= "----------------";	-- 0x014A
		when 000166 => D <= "----------------";	-- 0x014C
		when 000167 => D <= "----------------";	-- 0x014E
		when 000168 => D <= "----------------";	-- 0x0150
		when 000169 => D <= "----------------";	-- 0x0152
		when 000170 => D <= "----------------";	-- 0x0154
		when 000171 => D <= "----------------";	-- 0x0156
		when 000172 => D <= "----------------";	-- 0x0158
		when 000173 => D <= "----------------";	-- 0x015A
		when 000174 => D <= "----------------";	-- 0x015C
		when 000175 => D <= "----------------";	-- 0x015E
		when 000176 => D <= "----------------";	-- 0x0160
		when 000177 => D <= "----------------";	-- 0x0162
		when 000178 => D <= "----------------";	-- 0x0164
		when 000179 => D <= "----------------";	-- 0x0166
		when 000180 => D <= "----------------";	-- 0x0168
		when 000181 => D <= "----------------";	-- 0x016A
		when 000182 => D <= "----------------";	-- 0x016C
		when 000183 => D <= "----------------";	-- 0x016E
		when 000184 => D <= "----------------";	-- 0x0170
		when 000185 => D <= "----------------";	-- 0x0172
		when 000186 => D <= "----------------";	-- 0x0174
		when 000187 => D <= "----------------";	-- 0x0176
		when 000188 => D <= "----------------";	-- 0x0178
		when 000189 => D <= "----------------";	-- 0x017A
		when 000190 => D <= "----------------";	-- 0x017C
		when 000191 => D <= "----------------";	-- 0x017E
		when 000192 => D <= "----------------";	-- 0x0180
		when 000193 => D <= "----------------";	-- 0x0182
		when 000194 => D <= "----------------";	-- 0x0184
		when 000195 => D <= "----------------";	-- 0x0186
		when 000196 => D <= "----------------";	-- 0x0188
		when 000197 => D <= "----------------";	-- 0x018A
		when 000198 => D <= "----------------";	-- 0x018C
		when 000199 => D <= "----------------";	-- 0x018E
		when 000200 => D <= "----------------";	-- 0x0190
		when 000201 => D <= "----------------";	-- 0x0192
		when 000202 => D <= "----------------";	-- 0x0194
		when 000203 => D <= "----------------";	-- 0x0196
		when 000204 => D <= "----------------";	-- 0x0198
		when 000205 => D <= "----------------";	-- 0x019A
		when 000206 => D <= "----------------";	-- 0x019C
		when 000207 => D <= "----------------";	-- 0x019E
		when 000208 => D <= "----------------";	-- 0x01A0
		when 000209 => D <= "----------------";	-- 0x01A2
		when 000210 => D <= "----------------";	-- 0x01A4
		when 000211 => D <= "----------------";	-- 0x01A6
		when 000212 => D <= "----------------";	-- 0x01A8
		when 000213 => D <= "----------------";	-- 0x01AA
		when 000214 => D <= "----------------";	-- 0x01AC
		when 000215 => D <= "----------------";	-- 0x01AE
		when 000216 => D <= "----------------";	-- 0x01B0
		when 000217 => D <= "----------------";	-- 0x01B2
		when 000218 => D <= "----------------";	-- 0x01B4
		when 000219 => D <= "----------------";	-- 0x01B6
		when 000220 => D <= "----------------";	-- 0x01B8
		when 000221 => D <= "----------------";	-- 0x01BA
		when 000222 => D <= "----------------";	-- 0x01BC
		when 000223 => D <= "----------------";	-- 0x01BE
		when 000224 => D <= "----------------";	-- 0x01C0
		when 000225 => D <= "----------------";	-- 0x01C2
		when 000226 => D <= "----------------";	-- 0x01C4
		when 000227 => D <= "----------------";	-- 0x01C6
		when 000228 => D <= "----------------";	-- 0x01C8
		when 000229 => D <= "----------------";	-- 0x01CA
		when 000230 => D <= "----------------";	-- 0x01CC
		when 000231 => D <= "----------------";	-- 0x01CE
		when 000232 => D <= "----------------";	-- 0x01D0
		when 000233 => D <= "----------------";	-- 0x01D2
		when 000234 => D <= "----------------";	-- 0x01D4
		when 000235 => D <= "----------------";	-- 0x01D6
		when 000236 => D <= "----------------";	-- 0x01D8
		when 000237 => D <= "----------------";	-- 0x01DA
		when 000238 => D <= "----------------";	-- 0x01DC
		when 000239 => D <= "----------------";	-- 0x01DE
		when 000240 => D <= "----------------";	-- 0x01E0
		when 000241 => D <= "----------------";	-- 0x01E2
		when 000242 => D <= "----------------";	-- 0x01E4
		when 000243 => D <= "----------------";	-- 0x01E6
		when 000244 => D <= "----------------";	-- 0x01E8
		when 000245 => D <= "----------------";	-- 0x01EA
		when 000246 => D <= "----------------";	-- 0x01EC
		when 000247 => D <= "----------------";	-- 0x01EE
		when 000248 => D <= "----------------";	-- 0x01F0
		when 000249 => D <= "----------------";	-- 0x01F2
		when 000250 => D <= "----------------";	-- 0x01F4
		when 000251 => D <= "----------------";	-- 0x01F6
		when 000252 => D <= "----------------";	-- 0x01F8
		when 000253 => D <= "----------------";	-- 0x01FA
		when 000254 => D <= "----------------";	-- 0x01FC
		when 000255 => D <= "----------------";	-- 0x01FE
		when 000256 => D <= "----------------";	-- 0x0200
		when 000257 => D <= "----------------";	-- 0x0202
		when 000258 => D <= "----------------";	-- 0x0204
		when 000259 => D <= "----------------";	-- 0x0206
		when 000260 => D <= "----------------";	-- 0x0208
		when 000261 => D <= "----------------";	-- 0x020A
		when 000262 => D <= "----------------";	-- 0x020C
		when 000263 => D <= "----------------";	-- 0x020E
		when 000264 => D <= "----------------";	-- 0x0210
		when 000265 => D <= "----------------";	-- 0x0212
		when 000266 => D <= "----------------";	-- 0x0214
		when 000267 => D <= "----------------";	-- 0x0216
		when 000268 => D <= "----------------";	-- 0x0218
		when 000269 => D <= "----------------";	-- 0x021A
		when 000270 => D <= "----------------";	-- 0x021C
		when 000271 => D <= "----------------";	-- 0x021E
		when 000272 => D <= "----------------";	-- 0x0220
		when 000273 => D <= "----------------";	-- 0x0222
		when 000274 => D <= "----------------";	-- 0x0224
		when 000275 => D <= "----------------";	-- 0x0226
		when 000276 => D <= "----------------";	-- 0x0228
		when 000277 => D <= "----------------";	-- 0x022A
		when 000278 => D <= "----------------";	-- 0x022C
		when 000279 => D <= "----------------";	-- 0x022E
		when 000280 => D <= "----------------";	-- 0x0230
		when 000281 => D <= "----------------";	-- 0x0232
		when 000282 => D <= "----------------";	-- 0x0234
		when 000283 => D <= "----------------";	-- 0x0236
		when 000284 => D <= "----------------";	-- 0x0238
		when 000285 => D <= "----------------";	-- 0x023A
		when 000286 => D <= "----------------";	-- 0x023C
		when 000287 => D <= "----------------";	-- 0x023E
		when 000288 => D <= "----------------";	-- 0x0240
		when 000289 => D <= "----------------";	-- 0x0242
		when 000290 => D <= "----------------";	-- 0x0244
		when 000291 => D <= "----------------";	-- 0x0246
		when 000292 => D <= "----------------";	-- 0x0248
		when 000293 => D <= "----------------";	-- 0x024A
		when 000294 => D <= "----------------";	-- 0x024C
		when 000295 => D <= "----------------";	-- 0x024E
		when 000296 => D <= "----------------";	-- 0x0250
		when 000297 => D <= "----------------";	-- 0x0252
		when 000298 => D <= "----------------";	-- 0x0254
		when 000299 => D <= "----------------";	-- 0x0256
		when 000300 => D <= "----------------";	-- 0x0258
		when 000301 => D <= "----------------";	-- 0x025A
		when 000302 => D <= "----------------";	-- 0x025C
		when 000303 => D <= "----------------";	-- 0x025E
		when 000304 => D <= "----------------";	-- 0x0260
		when 000305 => D <= "----------------";	-- 0x0262
		when 000306 => D <= "----------------";	-- 0x0264
		when 000307 => D <= "----------------";	-- 0x0266
		when 000308 => D <= "----------------";	-- 0x0268
		when 000309 => D <= "----------------";	-- 0x026A
		when 000310 => D <= "----------------";	-- 0x026C
		when 000311 => D <= "----------------";	-- 0x026E
		when 000312 => D <= "----------------";	-- 0x0270
		when 000313 => D <= "----------------";	-- 0x0272
		when 000314 => D <= "----------------";	-- 0x0274
		when 000315 => D <= "----------------";	-- 0x0276
		when 000316 => D <= "----------------";	-- 0x0278
		when 000317 => D <= "----------------";	-- 0x027A
		when 000318 => D <= "----------------";	-- 0x027C
		when 000319 => D <= "----------------";	-- 0x027E
		when 000320 => D <= "----------------";	-- 0x0280
		when 000321 => D <= "----------------";	-- 0x0282
		when 000322 => D <= "----------------";	-- 0x0284
		when 000323 => D <= "----------------";	-- 0x0286
		when 000324 => D <= "----------------";	-- 0x0288
		when 000325 => D <= "----------------";	-- 0x028A
		when 000326 => D <= "----------------";	-- 0x028C
		when 000327 => D <= "----------------";	-- 0x028E
		when 000328 => D <= "----------------";	-- 0x0290
		when 000329 => D <= "----------------";	-- 0x0292
		when 000330 => D <= "----------------";	-- 0x0294
		when 000331 => D <= "----------------";	-- 0x0296
		when 000332 => D <= "----------------";	-- 0x0298
		when 000333 => D <= "----------------";	-- 0x029A
		when 000334 => D <= "----------------";	-- 0x029C
		when 000335 => D <= "----------------";	-- 0x029E
		when 000336 => D <= "----------------";	-- 0x02A0
		when 000337 => D <= "----------------";	-- 0x02A2
		when 000338 => D <= "----------------";	-- 0x02A4
		when 000339 => D <= "----------------";	-- 0x02A6
		when 000340 => D <= "----------------";	-- 0x02A8
		when 000341 => D <= "----------------";	-- 0x02AA
		when 000342 => D <= "----------------";	-- 0x02AC
		when 000343 => D <= "----------------";	-- 0x02AE
		when 000344 => D <= "----------------";	-- 0x02B0
		when 000345 => D <= "----------------";	-- 0x02B2
		when 000346 => D <= "----------------";	-- 0x02B4
		when 000347 => D <= "----------------";	-- 0x02B6
		when 000348 => D <= "----------------";	-- 0x02B8
		when 000349 => D <= "----------------";	-- 0x02BA
		when 000350 => D <= "----------------";	-- 0x02BC
		when 000351 => D <= "----------------";	-- 0x02BE
		when 000352 => D <= "----------------";	-- 0x02C0
		when 000353 => D <= "----------------";	-- 0x02C2
		when 000354 => D <= "----------------";	-- 0x02C4
		when 000355 => D <= "----------------";	-- 0x02C6
		when 000356 => D <= "----------------";	-- 0x02C8
		when 000357 => D <= "----------------";	-- 0x02CA
		when 000358 => D <= "----------------";	-- 0x02CC
		when 000359 => D <= "----------------";	-- 0x02CE
		when 000360 => D <= "----------------";	-- 0x02D0
		when 000361 => D <= "----------------";	-- 0x02D2
		when 000362 => D <= "----------------";	-- 0x02D4
		when 000363 => D <= "----------------";	-- 0x02D6
		when 000364 => D <= "----------------";	-- 0x02D8
		when 000365 => D <= "----------------";	-- 0x02DA
		when 000366 => D <= "----------------";	-- 0x02DC
		when 000367 => D <= "----------------";	-- 0x02DE
		when 000368 => D <= "----------------";	-- 0x02E0
		when 000369 => D <= "----------------";	-- 0x02E2
		when 000370 => D <= "----------------";	-- 0x02E4
		when 000371 => D <= "----------------";	-- 0x02E6
		when 000372 => D <= "----------------";	-- 0x02E8
		when 000373 => D <= "----------------";	-- 0x02EA
		when 000374 => D <= "----------------";	-- 0x02EC
		when 000375 => D <= "----------------";	-- 0x02EE
		when 000376 => D <= "----------------";	-- 0x02F0
		when 000377 => D <= "----------------";	-- 0x02F2
		when 000378 => D <= "----------------";	-- 0x02F4
		when 000379 => D <= "----------------";	-- 0x02F6
		when 000380 => D <= "----------------";	-- 0x02F8
		when 000381 => D <= "----------------";	-- 0x02FA
		when 000382 => D <= "----------------";	-- 0x02FC
		when 000383 => D <= "----------------";	-- 0x02FE
		when 000384 => D <= "----------------";	-- 0x0300
		when 000385 => D <= "----------------";	-- 0x0302
		when 000386 => D <= "----------------";	-- 0x0304
		when 000387 => D <= "----------------";	-- 0x0306
		when 000388 => D <= "----------------";	-- 0x0308
		when 000389 => D <= "----------------";	-- 0x030A
		when 000390 => D <= "----------------";	-- 0x030C
		when 000391 => D <= "----------------";	-- 0x030E
		when 000392 => D <= "----------------";	-- 0x0310
		when 000393 => D <= "----------------";	-- 0x0312
		when 000394 => D <= "----------------";	-- 0x0314
		when 000395 => D <= "----------------";	-- 0x0316
		when 000396 => D <= "----------------";	-- 0x0318
		when 000397 => D <= "----------------";	-- 0x031A
		when 000398 => D <= "----------------";	-- 0x031C
		when 000399 => D <= "----------------";	-- 0x031E
		when 000400 => D <= "----------------";	-- 0x0320
		when 000401 => D <= "----------------";	-- 0x0322
		when 000402 => D <= "----------------";	-- 0x0324
		when 000403 => D <= "----------------";	-- 0x0326
		when 000404 => D <= "----------------";	-- 0x0328
		when 000405 => D <= "----------------";	-- 0x032A
		when 000406 => D <= "----------------";	-- 0x032C
		when 000407 => D <= "----------------";	-- 0x032E
		when 000408 => D <= "----------------";	-- 0x0330
		when 000409 => D <= "----------------";	-- 0x0332
		when 000410 => D <= "----------------";	-- 0x0334
		when 000411 => D <= "----------------";	-- 0x0336
		when 000412 => D <= "----------------";	-- 0x0338
		when 000413 => D <= "----------------";	-- 0x033A
		when 000414 => D <= "----------------";	-- 0x033C
		when 000415 => D <= "----------------";	-- 0x033E
		when 000416 => D <= "----------------";	-- 0x0340
		when 000417 => D <= "----------------";	-- 0x0342
		when 000418 => D <= "----------------";	-- 0x0344
		when 000419 => D <= "----------------";	-- 0x0346
		when 000420 => D <= "----------------";	-- 0x0348
		when 000421 => D <= "----------------";	-- 0x034A
		when 000422 => D <= "----------------";	-- 0x034C
		when 000423 => D <= "----------------";	-- 0x034E
		when 000424 => D <= "----------------";	-- 0x0350
		when 000425 => D <= "----------------";	-- 0x0352
		when 000426 => D <= "----------------";	-- 0x0354
		when 000427 => D <= "----------------";	-- 0x0356
		when 000428 => D <= "----------------";	-- 0x0358
		when 000429 => D <= "----------------";	-- 0x035A
		when 000430 => D <= "----------------";	-- 0x035C
		when 000431 => D <= "----------------";	-- 0x035E
		when 000432 => D <= "----------------";	-- 0x0360
		when 000433 => D <= "----------------";	-- 0x0362
		when 000434 => D <= "----------------";	-- 0x0364
		when 000435 => D <= "----------------";	-- 0x0366
		when 000436 => D <= "----------------";	-- 0x0368
		when 000437 => D <= "----------------";	-- 0x036A
		when 000438 => D <= "----------------";	-- 0x036C
		when 000439 => D <= "----------------";	-- 0x036E
		when 000440 => D <= "----------------";	-- 0x0370
		when 000441 => D <= "----------------";	-- 0x0372
		when 000442 => D <= "----------------";	-- 0x0374
		when 000443 => D <= "----------------";	-- 0x0376
		when 000444 => D <= "----------------";	-- 0x0378
		when 000445 => D <= "----------------";	-- 0x037A
		when 000446 => D <= "----------------";	-- 0x037C
		when 000447 => D <= "----------------";	-- 0x037E
		when 000448 => D <= "----------------";	-- 0x0380
		when 000449 => D <= "----------------";	-- 0x0382
		when 000450 => D <= "----------------";	-- 0x0384
		when 000451 => D <= "----------------";	-- 0x0386
		when 000452 => D <= "----------------";	-- 0x0388
		when 000453 => D <= "----------------";	-- 0x038A
		when 000454 => D <= "----------------";	-- 0x038C
		when 000455 => D <= "----------------";	-- 0x038E
		when 000456 => D <= "----------------";	-- 0x0390
		when 000457 => D <= "----------------";	-- 0x0392
		when 000458 => D <= "----------------";	-- 0x0394
		when 000459 => D <= "----------------";	-- 0x0396
		when 000460 => D <= "----------------";	-- 0x0398
		when 000461 => D <= "----------------";	-- 0x039A
		when 000462 => D <= "----------------";	-- 0x039C
		when 000463 => D <= "----------------";	-- 0x039E
		when 000464 => D <= "----------------";	-- 0x03A0
		when 000465 => D <= "----------------";	-- 0x03A2
		when 000466 => D <= "----------------";	-- 0x03A4
		when 000467 => D <= "----------------";	-- 0x03A6
		when 000468 => D <= "----------------";	-- 0x03A8
		when 000469 => D <= "----------------";	-- 0x03AA
		when 000470 => D <= "----------------";	-- 0x03AC
		when 000471 => D <= "----------------";	-- 0x03AE
		when 000472 => D <= "----------------";	-- 0x03B0
		when 000473 => D <= "----------------";	-- 0x03B2
		when 000474 => D <= "----------------";	-- 0x03B4
		when 000475 => D <= "----------------";	-- 0x03B6
		when 000476 => D <= "----------------";	-- 0x03B8
		when 000477 => D <= "----------------";	-- 0x03BA
		when 000478 => D <= "----------------";	-- 0x03BC
		when 000479 => D <= "----------------";	-- 0x03BE
		when 000480 => D <= "----------------";	-- 0x03C0
		when 000481 => D <= "----------------";	-- 0x03C2
		when 000482 => D <= "----------------";	-- 0x03C4
		when 000483 => D <= "----------------";	-- 0x03C6
		when 000484 => D <= "----------------";	-- 0x03C8
		when 000485 => D <= "----------------";	-- 0x03CA
		when 000486 => D <= "----------------";	-- 0x03CC
		when 000487 => D <= "----------------";	-- 0x03CE
		when 000488 => D <= "----------------";	-- 0x03D0
		when 000489 => D <= "----------------";	-- 0x03D2
		when 000490 => D <= "----------------";	-- 0x03D4
		when 000491 => D <= "----------------";	-- 0x03D6
		when 000492 => D <= "----------------";	-- 0x03D8
		when 000493 => D <= "----------------";	-- 0x03DA
		when 000494 => D <= "----------------";	-- 0x03DC
		when 000495 => D <= "----------------";	-- 0x03DE
		when 000496 => D <= "----------------";	-- 0x03E0
		when 000497 => D <= "----------------";	-- 0x03E2
		when 000498 => D <= "----------------";	-- 0x03E4
		when 000499 => D <= "----------------";	-- 0x03E6
		when 000500 => D <= "----------------";	-- 0x03E8
		when 000501 => D <= "----------------";	-- 0x03EA
		when 000502 => D <= "----------------";	-- 0x03EC
		when 000503 => D <= "----------------";	-- 0x03EE
		when 000504 => D <= "----------------";	-- 0x03F0
		when 000505 => D <= "----------------";	-- 0x03F2
		when 000506 => D <= "----------------";	-- 0x03F4
		when 000507 => D <= "----------------";	-- 0x03F6
		when 000508 => D <= "----------------";	-- 0x03F8
		when 000509 => D <= "----------------";	-- 0x03FA
		when 000510 => D <= "----------------";	-- 0x03FC
		when 000511 => D <= "----------------";	-- 0x03FE
		when 000512 => D <= "0100000111111001";	-- 0x0400
		when 000513 => D <= "0000000000000001";	-- 0x0402
		when 000514 => D <= "0000000100000000";	-- 0x0404
		when 000515 => D <= "0100001000011000";	-- 0x0406
		when 000516 => D <= "1011000111111100";	-- 0x0408
		when 000517 => D <= "0000000000000001";	-- 0x040A
		when 000518 => D <= "0000000100100000";	-- 0x040C
		when 000519 => D <= "0110010111110110";	-- 0x040E
		when 000520 => D <= "0010001111000000";	-- 0x0410
		when 000521 => D <= "0000000000000001";	-- 0x0412
		when 000522 => D <= "0000000100001000";	-- 0x0414
		when 000523 => D <= "0010001111000001";	-- 0x0416
		when 000524 => D <= "0000000000000001";	-- 0x0418
		when 000525 => D <= "0000000100001100";	-- 0x041A
		when 000526 => D <= "0010001111111100";	-- 0x041C
		when 000527 => D <= "1111111111111111";	-- 0x041E
		when 000528 => D <= "1111111111111111";	-- 0x0420
		when 000529 => D <= "0000000000000001";	-- 0x0422
		when 000530 => D <= "0000000100000000";	-- 0x0424
		when 000531 => D <= "0010001111111100";	-- 0x0426
		when 000532 => D <= "0000000000000000";	-- 0x0428
		when 000533 => D <= "0000000000000000";	-- 0x042A
		when 000534 => D <= "0000000000000001";	-- 0x042C
		when 000535 => D <= "0000000100000100";	-- 0x042E
		when 000536 => D <= "0010001111111100";	-- 0x0430
		when 000537 => D <= "0000000000000001";	-- 0x0432
		when 000538 => D <= "0000000100100000";	-- 0x0434
		when 000539 => D <= "0000000000000001";	-- 0x0436
		when 000540 => D <= "0000000100010000";	-- 0x0438
		when 000541 => D <= "0010001111111100";	-- 0x043A
		when 000542 => D <= "0000000000000001";	-- 0x043C
		when 000543 => D <= "0011000000000000";	-- 0x043E
		when 000544 => D <= "0000000000000001";	-- 0x0440
		when 000545 => D <= "0000000100010100";	-- 0x0442
		when 000546 => D <= "0010111001111100";	-- 0x0444
		when 000547 => D <= "0000000000000001";	-- 0x0446
		when 000548 => D <= "0100000000000000";	-- 0x0448
		when 000549 => D <= "0100111010111001";	-- 0x044A
		when 000550 => D <= "0000000000000000";	-- 0x044C
		when 000551 => D <= "0000010010011100";	-- 0x044E
		when 000552 => D <= "0110000000010000";	-- 0x0450
		when 000553 => D <= "0100111001010110";	-- 0x0452
		when 000554 => D <= "0000000000000000";	-- 0x0454
		when 000555 => D <= "0010000000101110";	-- 0x0456
		when 000556 => D <= "0000000000001000";	-- 0x0458
		when 000557 => D <= "0100111001011110";	-- 0x045A
		when 000558 => D <= "1101111111111100";	-- 0x045C
		when 000559 => D <= "0000000000000000";	-- 0x045E
		when 000560 => D <= "0000000000001010";	-- 0x0460
		when 000561 => D <= "0100111001001111";	-- 0x0462
		when 000562 => D <= "0000000000000000";	-- 0x0464
		when 000563 => D <= "0110000010011000";	-- 0x0466
		when 000564 => D <= "0010000000101111";	-- 0x0468
		when 000565 => D <= "0000000000000100";	-- 0x046A
		when 000566 => D <= "0100111001001111";	-- 0x046C
		when 000567 => D <= "0000000000000001";	-- 0x046E
		when 000568 => D <= "0100111001110101";	-- 0x0470
		when 000569 => D <= "0100111001001111";	-- 0x0472
		when 000570 => D <= "0000000000000011";	-- 0x0474
		when 000571 => D <= "0100100010000000";	-- 0x0476
		when 000572 => D <= "0100100011000000";	-- 0x0478
		when 000573 => D <= "0100111001110101";	-- 0x047A
		when 000574 => D <= "0100111001001111";	-- 0x047C
		when 000575 => D <= "0000000000000100";	-- 0x047E
		when 000576 => D <= "0101011011000000";	-- 0x0480
		when 000577 => D <= "0100111001110101";	-- 0x0482
		when 000578 => D <= "0100111001001111";	-- 0x0484
		when 000579 => D <= "0000000000001001";	-- 0x0486
		when 000580 => D <= "0100111001110101";	-- 0x0488
		when 000581 => D <= "0100111111111001";	-- 0x048A
		when 000582 => D <= "0000000000000001";	-- 0x048C
		when 000583 => D <= "0100000000000000";	-- 0x048E
		when 000584 => D <= "0100000111111001";	-- 0x0490
		when 000585 => D <= "0000000000000000";	-- 0x0492
		when 000586 => D <= "0000010100101100";	-- 0x0494
		when 000587 => D <= "0100111001001111";	-- 0x0496
		when 000588 => D <= "0000000000000111";	-- 0x0498
		when 000589 => D <= "0110000011000110";	-- 0x049A
		when 000590 => D <= "0010111100001010";	-- 0x049C
		when 000591 => D <= "0100010111111001";	-- 0x049E
		when 000592 => D <= "0000000000000001";	-- 0x04A0
		when 000593 => D <= "0000000100011000";	-- 0x04A2
		when 000594 => D <= "0001001111111100";	-- 0x04A4
		when 000595 => D <= "0000000001100001";	-- 0x04A6
		when 000596 => D <= "0000000000000001";	-- 0x04A8
		when 000597 => D <= "0000000100011110";	-- 0x04AA
		when 000598 => D <= "0100001010010010";	-- 0x04AC
		when 000599 => D <= "0010000000010010";	-- 0x04AE
		when 000600 => D <= "0110011000000000";	-- 0x04B0
		when 000601 => D <= "0000000001110110";	-- 0x04B2
		when 000602 => D <= "0010000001111001";	-- 0x04B4
		when 000603 => D <= "0000000000000000";	-- 0x04B6
		when 000604 => D <= "0000010101010110";	-- 0x04B8
		when 000605 => D <= "0001000000010000";	-- 0x04BA
		when 000606 => D <= "1100000000111100";	-- 0x04BC
		when 000607 => D <= "0000000000001000";	-- 0x04BE
		when 000608 => D <= "0110011100010100";	-- 0x04C0
		when 000609 => D <= "0010000001111001";	-- 0x04C2
		when 000610 => D <= "0000000000000000";	-- 0x04C4
		when 000611 => D <= "0000010101010010";	-- 0x04C6
		when 000612 => D <= "0001000010111001";	-- 0x04C8
		when 000613 => D <= "0000000000000001";	-- 0x04CA
		when 000614 => D <= "0000000100011110";	-- 0x04CC
		when 000615 => D <= "0101001000111001";	-- 0x04CE
		when 000616 => D <= "0000000000000001";	-- 0x04D0
		when 000617 => D <= "0000000100011110";	-- 0x04D2
		when 000618 => D <= "0110000000111100";	-- 0x04D4
		when 000619 => D <= "0010000001111001";	-- 0x04D6
		when 000620 => D <= "0000000000000000";	-- 0x04D8
		when 000621 => D <= "0000010101010110";	-- 0x04DA
		when 000622 => D <= "0001000000010000";	-- 0x04DC
		when 000623 => D <= "1100000000111100";	-- 0x04DE
		when 000624 => D <= "0000000000000001";	-- 0x04E0
		when 000625 => D <= "0110011100101110";	-- 0x04E2
		when 000626 => D <= "0010000001111001";	-- 0x04E4
		when 000627 => D <= "0000000000000000";	-- 0x04E6
		when 000628 => D <= "0000010101010010";	-- 0x04E8
		when 000629 => D <= "0001001111010000";	-- 0x04EA
		when 000630 => D <= "0000000000000001";	-- 0x04EC
		when 000631 => D <= "0000000100011100";	-- 0x04EE
		when 000632 => D <= "0001000000111001";	-- 0x04F0
		when 000633 => D <= "0000000000000001";	-- 0x04F2
		when 000634 => D <= "0000000100011100";	-- 0x04F4
		when 000635 => D <= "0100100010000000";	-- 0x04F6
		when 000636 => D <= "0100100011000000";	-- 0x04F8
		when 000637 => D <= "0100000111111001";	-- 0x04FA
		when 000638 => D <= "0000000000000000";	-- 0x04FC
		when 000639 => D <= "0000010101010000";	-- 0x04FE
		when 000640 => D <= "1011000010001000";	-- 0x0500
		when 000641 => D <= "0110011000001110";	-- 0x0502
		when 000642 => D <= "0001001111111100";	-- 0x0504
		when 000643 => D <= "0000000001100001";	-- 0x0506
		when 000644 => D <= "0000000000000001";	-- 0x0508
		when 000645 => D <= "0000000100011110";	-- 0x050A
		when 000646 => D <= "0010010010111100";	-- 0x050C
		when 000647 => D <= "0000000000000000";	-- 0x050E
		when 000648 => D <= "0000000000000001";	-- 0x0510
		when 000649 => D <= "0001000000111001";	-- 0x0512
		when 000650 => D <= "0000000000000001";	-- 0x0514
		when 000651 => D <= "0000000100011110";	-- 0x0516
		when 000652 => D <= "0000110000000000";	-- 0x0518
		when 000653 => D <= "0000000001111010";	-- 0x051A
		when 000654 => D <= "0110111100001000";	-- 0x051C
		when 000655 => D <= "0001001111111100";	-- 0x051E
		when 000656 => D <= "0000000001100001";	-- 0x0520
		when 000657 => D <= "0000000000000001";	-- 0x0522
		when 000658 => D <= "0000000100011110";	-- 0x0524
		when 000659 => D <= "0110000010000110";	-- 0x0526
		when 000660 => D <= "0010010001011111";	-- 0x0528
		when 000661 => D <= "0100111001110101";	-- 0x052A
		when 000662 => D <= "0101001101110100";	-- 0x052C
		when 000663 => D <= "0110000101100011";	-- 0x052E
		when 000664 => D <= "0110101100100000";	-- 0x0530
		when 000665 => D <= "0110111101110110";	-- 0x0532
		when 000666 => D <= "0110010101110010";	-- 0x0534
		when 000667 => D <= "0110011001101100";	-- 0x0536
		when 000668 => D <= "0110111101110111";	-- 0x0538
		when 000669 => D <= "0010000100001010";	-- 0x053A
		when 000670 => D <= "0000110101010000";	-- 0x053C
		when 000671 => D <= "0111001001101111";	-- 0x053E
		when 000672 => D <= "0110011101110010";	-- 0x0540
		when 000673 => D <= "0110000101101101";	-- 0x0542
		when 000674 => D <= "0010000001100001";	-- 0x0544
		when 000675 => D <= "0110001001101111";	-- 0x0546
		when 000676 => D <= "0111001001110100";	-- 0x0548
		when 000677 => D <= "0110010101100100";	-- 0x054A
		when 000678 => D <= "0000101000001101";	-- 0x054C
		when 000679 => D <= "0000000000000000";	-- 0x054E
		when 000680 => D <= "0111001100000000";	-- 0x0550
		when 000681 => D <= "0000000000001000";	-- 0x0552
		when 000682 => D <= "0000000000000000";	-- 0x0554
		when 000683 => D <= "0000000000001000";	-- 0x0556
		when 000684 => D <= "0000000000000010";	-- 0x0558
		when others => D <= "----------------";
		end case;
	end process;
end;
