-- This file was generated with hex2rom written by Daniel Wallner

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
	port(
		A	: in std_logic_vector(11 downto 0);
		D	: out std_logic_vector(15 downto 0)
	);
end rom;

architecture rtl of rom is
begin
	process (A)
	begin
		case to_integer(unsigned(A)) is
		when 000000 => D <= "0000000000000001";	-- 0x0000
		when 000001 => D <= "0111111111111110";	-- 0x0002
		when 000002 => D <= "0000000000000000";	-- 0x0004
		when 000003 => D <= "0000000100000000";	-- 0x0006
		when 000004 => D <= "0000000000000000";	-- 0x0008
		when 000005 => D <= "0000000000000000";	-- 0x000A
		when 000006 => D <= "0000000000000000";	-- 0x000C
		when 000007 => D <= "0000000110000000";	-- 0x000E
		when 000008 => D <= "0000000000000000";	-- 0x0010
		when 000009 => D <= "0000000110000100";	-- 0x0012
		when 000010 => D <= "----------------";	-- 0x0014
		when 000011 => D <= "----------------";	-- 0x0016
		when 000012 => D <= "----------------";	-- 0x0018
		when 000013 => D <= "----------------";	-- 0x001A
		when 000014 => D <= "----------------";	-- 0x001C
		when 000015 => D <= "----------------";	-- 0x001E
		when 000016 => D <= "----------------";	-- 0x0020
		when 000017 => D <= "----------------";	-- 0x0022
		when 000018 => D <= "----------------";	-- 0x0024
		when 000019 => D <= "----------------";	-- 0x0026
		when 000020 => D <= "----------------";	-- 0x0028
		when 000021 => D <= "----------------";	-- 0x002A
		when 000022 => D <= "----------------";	-- 0x002C
		when 000023 => D <= "----------------";	-- 0x002E
		when 000024 => D <= "----------------";	-- 0x0030
		when 000025 => D <= "----------------";	-- 0x0032
		when 000026 => D <= "----------------";	-- 0x0034
		when 000027 => D <= "----------------";	-- 0x0036
		when 000028 => D <= "----------------";	-- 0x0038
		when 000029 => D <= "----------------";	-- 0x003A
		when 000030 => D <= "----------------";	-- 0x003C
		when 000031 => D <= "----------------";	-- 0x003E
		when 000032 => D <= "----------------";	-- 0x0040
		when 000033 => D <= "----------------";	-- 0x0042
		when 000034 => D <= "----------------";	-- 0x0044
		when 000035 => D <= "----------------";	-- 0x0046
		when 000036 => D <= "----------------";	-- 0x0048
		when 000037 => D <= "----------------";	-- 0x004A
		when 000038 => D <= "----------------";	-- 0x004C
		when 000039 => D <= "----------------";	-- 0x004E
		when 000040 => D <= "----------------";	-- 0x0050
		when 000041 => D <= "----------------";	-- 0x0052
		when 000042 => D <= "----------------";	-- 0x0054
		when 000043 => D <= "----------------";	-- 0x0056
		when 000044 => D <= "----------------";	-- 0x0058
		when 000045 => D <= "----------------";	-- 0x005A
		when 000046 => D <= "----------------";	-- 0x005C
		when 000047 => D <= "----------------";	-- 0x005E
		when 000048 => D <= "----------------";	-- 0x0060
		when 000049 => D <= "----------------";	-- 0x0062
		when 000050 => D <= "----------------";	-- 0x0064
		when 000051 => D <= "----------------";	-- 0x0066
		when 000052 => D <= "----------------";	-- 0x0068
		when 000053 => D <= "----------------";	-- 0x006A
		when 000054 => D <= "----------------";	-- 0x006C
		when 000055 => D <= "----------------";	-- 0x006E
		when 000056 => D <= "----------------";	-- 0x0070
		when 000057 => D <= "----------------";	-- 0x0072
		when 000058 => D <= "----------------";	-- 0x0074
		when 000059 => D <= "----------------";	-- 0x0076
		when 000060 => D <= "----------------";	-- 0x0078
		when 000061 => D <= "----------------";	-- 0x007A
		when 000062 => D <= "----------------";	-- 0x007C
		when 000063 => D <= "----------------";	-- 0x007E
		when 000064 => D <= "----------------";	-- 0x0080
		when 000065 => D <= "----------------";	-- 0x0082
		when 000066 => D <= "----------------";	-- 0x0084
		when 000067 => D <= "----------------";	-- 0x0086
		when 000068 => D <= "----------------";	-- 0x0088
		when 000069 => D <= "----------------";	-- 0x008A
		when 000070 => D <= "----------------";	-- 0x008C
		when 000071 => D <= "----------------";	-- 0x008E
		when 000072 => D <= "----------------";	-- 0x0090
		when 000073 => D <= "----------------";	-- 0x0092
		when 000074 => D <= "----------------";	-- 0x0094
		when 000075 => D <= "----------------";	-- 0x0096
		when 000076 => D <= "----------------";	-- 0x0098
		when 000077 => D <= "----------------";	-- 0x009A
		when 000078 => D <= "----------------";	-- 0x009C
		when 000079 => D <= "----------------";	-- 0x009E
		when 000080 => D <= "----------------";	-- 0x00A0
		when 000081 => D <= "----------------";	-- 0x00A2
		when 000082 => D <= "----------------";	-- 0x00A4
		when 000083 => D <= "----------------";	-- 0x00A6
		when 000084 => D <= "----------------";	-- 0x00A8
		when 000085 => D <= "----------------";	-- 0x00AA
		when 000086 => D <= "----------------";	-- 0x00AC
		when 000087 => D <= "----------------";	-- 0x00AE
		when 000088 => D <= "----------------";	-- 0x00B0
		when 000089 => D <= "----------------";	-- 0x00B2
		when 000090 => D <= "----------------";	-- 0x00B4
		when 000091 => D <= "----------------";	-- 0x00B6
		when 000092 => D <= "----------------";	-- 0x00B8
		when 000093 => D <= "----------------";	-- 0x00BA
		when 000094 => D <= "----------------";	-- 0x00BC
		when 000095 => D <= "----------------";	-- 0x00BE
		when 000096 => D <= "----------------";	-- 0x00C0
		when 000097 => D <= "----------------";	-- 0x00C2
		when 000098 => D <= "----------------";	-- 0x00C4
		when 000099 => D <= "----------------";	-- 0x00C6
		when 000100 => D <= "----------------";	-- 0x00C8
		when 000101 => D <= "----------------";	-- 0x00CA
		when 000102 => D <= "----------------";	-- 0x00CC
		when 000103 => D <= "----------------";	-- 0x00CE
		when 000104 => D <= "----------------";	-- 0x00D0
		when 000105 => D <= "----------------";	-- 0x00D2
		when 000106 => D <= "----------------";	-- 0x00D4
		when 000107 => D <= "----------------";	-- 0x00D6
		when 000108 => D <= "----------------";	-- 0x00D8
		when 000109 => D <= "----------------";	-- 0x00DA
		when 000110 => D <= "----------------";	-- 0x00DC
		when 000111 => D <= "----------------";	-- 0x00DE
		when 000112 => D <= "----------------";	-- 0x00E0
		when 000113 => D <= "----------------";	-- 0x00E2
		when 000114 => D <= "----------------";	-- 0x00E4
		when 000115 => D <= "----------------";	-- 0x00E6
		when 000116 => D <= "----------------";	-- 0x00E8
		when 000117 => D <= "----------------";	-- 0x00EA
		when 000118 => D <= "----------------";	-- 0x00EC
		when 000119 => D <= "----------------";	-- 0x00EE
		when 000120 => D <= "----------------";	-- 0x00F0
		when 000121 => D <= "----------------";	-- 0x00F2
		when 000122 => D <= "----------------";	-- 0x00F4
		when 000123 => D <= "----------------";	-- 0x00F6
		when 000124 => D <= "----------------";	-- 0x00F8
		when 000125 => D <= "----------------";	-- 0x00FA
		when 000126 => D <= "----------------";	-- 0x00FC
		when 000127 => D <= "----------------";	-- 0x00FE
		when 000128 => D <= "0010111001111000";	-- 0x0100
		when 000129 => D <= "0000000000000000";	-- 0x0102
		when 000130 => D <= "0011111100111100";	-- 0x0104
		when 000131 => D <= "0101010110001000";	-- 0x0106
		when 000132 => D <= "0011000000011111";	-- 0x0108
		when 000133 => D <= "0010101001111100";	-- 0x010A
		when 000134 => D <= "0000000000000001";	-- 0x010C
		when 000135 => D <= "0000000000000000";	-- 0x010E
		when 000136 => D <= "0010001111111100";	-- 0x0110
		when 000137 => D <= "0001001000110100";	-- 0x0112
		when 000138 => D <= "0101011001111000";	-- 0x0114
		when 000139 => D <= "0000000000000001";	-- 0x0116
		when 000140 => D <= "0000000000000000";	-- 0x0118
		when 000141 => D <= "0010101011111100";	-- 0x011A
		when 000142 => D <= "1011000000001011";	-- 0x011C
		when 000143 => D <= "1111000000001101";	-- 0x011E
		when 000144 => D <= "0010101010111100";	-- 0x0120
		when 000145 => D <= "1101111010101101";	-- 0x0122
		when 000146 => D <= "1011111011101111";	-- 0x0124
		when 000147 => D <= "0001001111111100";	-- 0x0126
		when 000148 => D <= "0000000000001010";	-- 0x0128
		when 000149 => D <= "0000000000000001";	-- 0x012A
		when 000150 => D <= "0000000100000000";	-- 0x012C
		when 000151 => D <= "0001001111111100";	-- 0x012E
		when 000152 => D <= "0000000000001011";	-- 0x0130
		when 000153 => D <= "0000000000000001";	-- 0x0132
		when 000154 => D <= "0000000100000001";	-- 0x0134
		when 000155 => D <= "0001001111111100";	-- 0x0136
		when 000156 => D <= "0000000000001100";	-- 0x0138
		when 000157 => D <= "0000000000000001";	-- 0x013A
		when 000158 => D <= "0000000100000010";	-- 0x013C
		when 000159 => D <= "0001001111111100";	-- 0x013E
		when 000160 => D <= "0000000000001101";	-- 0x0140
		when 000161 => D <= "0000000000000001";	-- 0x0142
		when 000162 => D <= "0000000100000011";	-- 0x0144
		when 000163 => D <= "0011011000111001";	-- 0x0146
		when 000164 => D <= "0000000000000001";	-- 0x0148
		when 000165 => D <= "0000000100000000";	-- 0x014A
		when 000166 => D <= "0010011000111001";	-- 0x014C
		when 000167 => D <= "0000000000000001";	-- 0x014E
		when 000168 => D <= "0000000100000000";	-- 0x0150
		when 000169 => D <= "0010001111000011";	-- 0x0152
		when 000170 => D <= "0000000000000001";	-- 0x0154
		when 000171 => D <= "0000000000100000";	-- 0x0156
		when 000172 => D <= "0001011000111100";	-- 0x0158
		when 000173 => D <= "0000000001000001";	-- 0x015A
		when 000174 => D <= "0010011001111100";	-- 0x015C
		when 000175 => D <= "0000000000001000";	-- 0x015E
		when 000176 => D <= "0000000000000000";	-- 0x0160
		when 000177 => D <= "0010100001111100";	-- 0x0162
		when 000178 => D <= "0000000000001000";	-- 0x0164
		when 000179 => D <= "0000000000000010";	-- 0x0166
		when 000180 => D <= "0001011010000011";	-- 0x0168
		when 000181 => D <= "0010101000010101";	-- 0x016A
		when 000182 => D <= "0001100000010100";	-- 0x016C
		when 000183 => D <= "0000100000000100";	-- 0x016E
		when 000184 => D <= "0000000000010000";	-- 0x0170
		when 000185 => D <= "0110011111111000";	-- 0x0172
		when 000186 => D <= "0100111001110001";	-- 0x0174
		when 000187 => D <= "0100111001110001";	-- 0x0176
		when 000188 => D <= "0100111001110001";	-- 0x0178
		when 000189 => D <= "0100111001110001";	-- 0x017A
		when 000190 => D <= "0100111011111000";	-- 0x017C
		when 000191 => D <= "0000000100000000";	-- 0x017E
		when 000192 => D <= "0100111011111000";	-- 0x0180
		when 000193 => D <= "0000000110000000";	-- 0x0182
		when 000194 => D <= "0100111011111000";	-- 0x0184
		when 000195 => D <= "0000000110000100";	-- 0x0186
		when others => D <= "----------------";
		end case;
	end process;
end;
