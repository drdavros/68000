-- This file was generated with hex2rom written by Daniel Wallner

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom is
	port(
		A	: in std_logic_vector(11 downto 0);
		D	: out std_logic_vector(15 downto 0)
	);
end rom;

architecture rtl of rom is
begin
	process (A)
	begin
		case to_integer(unsigned(A)) is
		when 000000 => D <= "0000000000000001";	-- 0x0000
		when 000001 => D <= "0011111111111110";	-- 0x0002
		when 000002 => D <= "0000000000000000";	-- 0x0004
		when 000003 => D <= "0000000100100000";	-- 0x0006
		when 000004 => D <= "----------------";	-- 0x0008
		when 000005 => D <= "----------------";	-- 0x000A
		when 000006 => D <= "----------------";	-- 0x000C
		when 000007 => D <= "----------------";	-- 0x000E
		when 000008 => D <= "----------------";	-- 0x0010
		when 000009 => D <= "----------------";	-- 0x0012
		when 000010 => D <= "----------------";	-- 0x0014
		when 000011 => D <= "----------------";	-- 0x0016
		when 000012 => D <= "----------------";	-- 0x0018
		when 000013 => D <= "----------------";	-- 0x001A
		when 000014 => D <= "----------------";	-- 0x001C
		when 000015 => D <= "----------------";	-- 0x001E
		when 000016 => D <= "----------------";	-- 0x0020
		when 000017 => D <= "----------------";	-- 0x0022
		when 000018 => D <= "----------------";	-- 0x0024
		when 000019 => D <= "----------------";	-- 0x0026
		when 000020 => D <= "----------------";	-- 0x0028
		when 000021 => D <= "----------------";	-- 0x002A
		when 000022 => D <= "----------------";	-- 0x002C
		when 000023 => D <= "----------------";	-- 0x002E
		when 000024 => D <= "----------------";	-- 0x0030
		when 000025 => D <= "----------------";	-- 0x0032
		when 000026 => D <= "----------------";	-- 0x0034
		when 000027 => D <= "----------------";	-- 0x0036
		when 000028 => D <= "----------------";	-- 0x0038
		when 000029 => D <= "----------------";	-- 0x003A
		when 000030 => D <= "----------------";	-- 0x003C
		when 000031 => D <= "----------------";	-- 0x003E
		when 000032 => D <= "----------------";	-- 0x0040
		when 000033 => D <= "----------------";	-- 0x0042
		when 000034 => D <= "----------------";	-- 0x0044
		when 000035 => D <= "----------------";	-- 0x0046
		when 000036 => D <= "----------------";	-- 0x0048
		when 000037 => D <= "----------------";	-- 0x004A
		when 000038 => D <= "----------------";	-- 0x004C
		when 000039 => D <= "----------------";	-- 0x004E
		when 000040 => D <= "----------------";	-- 0x0050
		when 000041 => D <= "----------------";	-- 0x0052
		when 000042 => D <= "----------------";	-- 0x0054
		when 000043 => D <= "----------------";	-- 0x0056
		when 000044 => D <= "----------------";	-- 0x0058
		when 000045 => D <= "----------------";	-- 0x005A
		when 000046 => D <= "----------------";	-- 0x005C
		when 000047 => D <= "----------------";	-- 0x005E
		when 000048 => D <= "----------------";	-- 0x0060
		when 000049 => D <= "----------------";	-- 0x0062
		when 000050 => D <= "----------------";	-- 0x0064
		when 000051 => D <= "----------------";	-- 0x0066
		when 000052 => D <= "----------------";	-- 0x0068
		when 000053 => D <= "----------------";	-- 0x006A
		when 000054 => D <= "----------------";	-- 0x006C
		when 000055 => D <= "----------------";	-- 0x006E
		when 000056 => D <= "----------------";	-- 0x0070
		when 000057 => D <= "----------------";	-- 0x0072
		when 000058 => D <= "----------------";	-- 0x0074
		when 000059 => D <= "----------------";	-- 0x0076
		when 000060 => D <= "----------------";	-- 0x0078
		when 000061 => D <= "----------------";	-- 0x007A
		when 000062 => D <= "----------------";	-- 0x007C
		when 000063 => D <= "----------------";	-- 0x007E
		when 000064 => D <= "----------------";	-- 0x0080
		when 000065 => D <= "----------------";	-- 0x0082
		when 000066 => D <= "----------------";	-- 0x0084
		when 000067 => D <= "----------------";	-- 0x0086
		when 000068 => D <= "----------------";	-- 0x0088
		when 000069 => D <= "----------------";	-- 0x008A
		when 000070 => D <= "----------------";	-- 0x008C
		when 000071 => D <= "----------------";	-- 0x008E
		when 000072 => D <= "----------------";	-- 0x0090
		when 000073 => D <= "----------------";	-- 0x0092
		when 000074 => D <= "----------------";	-- 0x0094
		when 000075 => D <= "----------------";	-- 0x0096
		when 000076 => D <= "----------------";	-- 0x0098
		when 000077 => D <= "----------------";	-- 0x009A
		when 000078 => D <= "----------------";	-- 0x009C
		when 000079 => D <= "----------------";	-- 0x009E
		when 000080 => D <= "----------------";	-- 0x00A0
		when 000081 => D <= "----------------";	-- 0x00A2
		when 000082 => D <= "----------------";	-- 0x00A4
		when 000083 => D <= "----------------";	-- 0x00A6
		when 000084 => D <= "----------------";	-- 0x00A8
		when 000085 => D <= "----------------";	-- 0x00AA
		when 000086 => D <= "----------------";	-- 0x00AC
		when 000087 => D <= "----------------";	-- 0x00AE
		when 000088 => D <= "----------------";	-- 0x00B0
		when 000089 => D <= "----------------";	-- 0x00B2
		when 000090 => D <= "----------------";	-- 0x00B4
		when 000091 => D <= "----------------";	-- 0x00B6
		when 000092 => D <= "----------------";	-- 0x00B8
		when 000093 => D <= "----------------";	-- 0x00BA
		when 000094 => D <= "----------------";	-- 0x00BC
		when 000095 => D <= "----------------";	-- 0x00BE
		when 000096 => D <= "----------------";	-- 0x00C0
		when 000097 => D <= "----------------";	-- 0x00C2
		when 000098 => D <= "----------------";	-- 0x00C4
		when 000099 => D <= "----------------";	-- 0x00C6
		when 000100 => D <= "----------------";	-- 0x00C8
		when 000101 => D <= "----------------";	-- 0x00CA
		when 000102 => D <= "----------------";	-- 0x00CC
		when 000103 => D <= "----------------";	-- 0x00CE
		when 000104 => D <= "----------------";	-- 0x00D0
		when 000105 => D <= "----------------";	-- 0x00D2
		when 000106 => D <= "----------------";	-- 0x00D4
		when 000107 => D <= "----------------";	-- 0x00D6
		when 000108 => D <= "----------------";	-- 0x00D8
		when 000109 => D <= "----------------";	-- 0x00DA
		when 000110 => D <= "----------------";	-- 0x00DC
		when 000111 => D <= "----------------";	-- 0x00DE
		when 000112 => D <= "----------------";	-- 0x00E0
		when 000113 => D <= "----------------";	-- 0x00E2
		when 000114 => D <= "----------------";	-- 0x00E4
		when 000115 => D <= "----------------";	-- 0x00E6
		when 000116 => D <= "----------------";	-- 0x00E8
		when 000117 => D <= "----------------";	-- 0x00EA
		when 000118 => D <= "----------------";	-- 0x00EC
		when 000119 => D <= "----------------";	-- 0x00EE
		when 000120 => D <= "----------------";	-- 0x00F0
		when 000121 => D <= "----------------";	-- 0x00F2
		when 000122 => D <= "----------------";	-- 0x00F4
		when 000123 => D <= "----------------";	-- 0x00F6
		when 000124 => D <= "----------------";	-- 0x00F8
		when 000125 => D <= "----------------";	-- 0x00FA
		when 000126 => D <= "----------------";	-- 0x00FC
		when 000127 => D <= "----------------";	-- 0x00FE
		when 000128 => D <= "0000000000000001";	-- 0x0100
		when 000129 => D <= "0000000010000000";	-- 0x0102
		when 000130 => D <= "0110000000000000";	-- 0x0104
		when 000131 => D <= "0000000000100100";	-- 0x0106
		when 000132 => D <= "0110000000000000";	-- 0x0108
		when 000133 => D <= "0000000001010010";	-- 0x010A
		when 000134 => D <= "0110000000000000";	-- 0x010C
		when 000135 => D <= "0000110010101100";	-- 0x010E
		when 000136 => D <= "0110000000000000";	-- 0x0110
		when 000137 => D <= "0000110010111010";	-- 0x0112
		when 000138 => D <= "0110000000000000";	-- 0x0114
		when 000139 => D <= "0000110011001110";	-- 0x0116
		when 000140 => D <= "0110000000000000";	-- 0x0118
		when 000141 => D <= "0000110011011100";	-- 0x011A
		when 000142 => D <= "0110000000000000";	-- 0x011C
		when 000143 => D <= "0000110011110000";	-- 0x011E
		when 000144 => D <= "0010001111111100";	-- 0x0120
		when 000145 => D <= "0000000000000000";	-- 0x0122
		when 000146 => D <= "0000000100000100";	-- 0x0124
		when 000147 => D <= "0000000000000001";	-- 0x0126
		when 000148 => D <= "0000000000000000";	-- 0x0128
		when 000149 => D <= "0010111001111000";	-- 0x012A
		when 000150 => D <= "0000000000000000";	-- 0x012C
		when 000151 => D <= "0100110111111001";	-- 0x012E
		when 000152 => D <= "0000000000000000";	-- 0x0130
		when 000153 => D <= "0000111000010100";	-- 0x0132
		when 000154 => D <= "0110000100000000";	-- 0x0134
		when 000155 => D <= "0000110001110110";	-- 0x0136
		when 000156 => D <= "0010001111111000";	-- 0x0138
		when 000157 => D <= "0000000100000000";	-- 0x013A
		when 000158 => D <= "0000000000000001";	-- 0x013C
		when 000159 => D <= "0000000000100100";	-- 0x013E
		when 000160 => D <= "0010000000111000";	-- 0x0140
		when 000161 => D <= "0000000000000000";	-- 0x0142
		when 000162 => D <= "0000010010000000";	-- 0x0144
		when 000163 => D <= "0000000000000000";	-- 0x0146
		when 000164 => D <= "0000100000000000";	-- 0x0148
		when 000165 => D <= "0010001111000000";	-- 0x014A
		when 000166 => D <= "0000000000000001";	-- 0x014C
		when 000167 => D <= "0000000000101100";	-- 0x014E
		when 000168 => D <= "0000010010000000";	-- 0x0150
		when 000169 => D <= "0000000000000000";	-- 0x0152
		when 000170 => D <= "0000000001101100";	-- 0x0154
		when 000171 => D <= "0010001111000000";	-- 0x0156
		when 000172 => D <= "0000000000000001";	-- 0x0158
		when 000173 => D <= "0000000000101000";	-- 0x015A
		when 000174 => D <= "0100001010000000";	-- 0x015C
		when 000175 => D <= "0010001111000000";	-- 0x015E
		when 000176 => D <= "0000000000000001";	-- 0x0160
		when 000177 => D <= "0000000000010000";	-- 0x0162
		when 000178 => D <= "0010001111000000";	-- 0x0164
		when 000179 => D <= "0000000000000001";	-- 0x0166
		when 000180 => D <= "0000000000001000";	-- 0x0168
		when 000181 => D <= "0010001111000000";	-- 0x016A
		when 000182 => D <= "0000000000000001";	-- 0x016C
		when 000183 => D <= "0000000000000100";	-- 0x016E
		when 000184 => D <= "0010111001111000";	-- 0x0170
		when 000185 => D <= "0000000000000000";	-- 0x0172
		when 000186 => D <= "0100110111111001";	-- 0x0174
		when 000187 => D <= "0000000000000000";	-- 0x0176
		when 000188 => D <= "0000111000111010";	-- 0x0178
		when 000189 => D <= "0110000100000000";	-- 0x017A
		when 000190 => D <= "0000110000110000";	-- 0x017C
		when 000191 => D <= "0001000000111100";	-- 0x017E
		when 000192 => D <= "0000000000111110";	-- 0x0180
		when 000193 => D <= "0110000100000000";	-- 0x0182
		when 000194 => D <= "0000100100000010";	-- 0x0184
		when 000195 => D <= "0110000100000000";	-- 0x0186
		when 000196 => D <= "0000101110101110";	-- 0x0188
		when 000197 => D <= "0010100001001000";	-- 0x018A
		when 000198 => D <= "0100000111111001";	-- 0x018C
		when 000199 => D <= "0000000000000001";	-- 0x018E
		when 000200 => D <= "0000000000110000";	-- 0x0190
		when 000201 => D <= "0110000100000000";	-- 0x0192
		when 000202 => D <= "0000101101011000";	-- 0x0194
		when 000203 => D <= "0110000100000000";	-- 0x0196
		when 000204 => D <= "0000101110010000";	-- 0x0198
		when 000205 => D <= "0100101001000001";	-- 0x019A
		when 000206 => D <= "0110011100000000";	-- 0x019C
		when 000207 => D <= "0000000101101110";	-- 0x019E
		when 000208 => D <= "1011001010111100";	-- 0x01A0
		when 000209 => D <= "0000000000000000";	-- 0x01A2
		when 000210 => D <= "1111111111111111";	-- 0x01A4
		when 000211 => D <= "0110010000000000";	-- 0x01A6
		when 000212 => D <= "0000100011010100";	-- 0x01A8
		when 000213 => D <= "0001000100000001";	-- 0x01AA
		when 000214 => D <= "1110000001011001";	-- 0x01AC
		when 000215 => D <= "0001000100000001";	-- 0x01AE
		when 000216 => D <= "1110000101011001";	-- 0x01B0
		when 000217 => D <= "0110000100000000";	-- 0x01B2
		when 000218 => D <= "0000100110000000";	-- 0x01B4
		when 000219 => D <= "0010101001001001";	-- 0x01B6
		when 000220 => D <= "0110011000000000";	-- 0x01B8
		when 000221 => D <= "0000000000011000";	-- 0x01BA
		when 000222 => D <= "0110000100000000";	-- 0x01BC
		when 000223 => D <= "0000100110100010";	-- 0x01BE
		when 000224 => D <= "0010010001001101";	-- 0x01C0
		when 000225 => D <= "0010011001111001";	-- 0x01C2
		when 000226 => D <= "0000000000000001";	-- 0x01C4
		when 000227 => D <= "0000000000100100";	-- 0x01C6
		when 000228 => D <= "0110000100000000";	-- 0x01C8
		when 000229 => D <= "0000100110100000";	-- 0x01CA
		when 000230 => D <= "0010001111001010";	-- 0x01CC
		when 000231 => D <= "0000000000000001";	-- 0x01CE
		when 000232 => D <= "0000000000100100";	-- 0x01D0
		when 000233 => D <= "0010000000001100";	-- 0x01D2
		when 000234 => D <= "1001000010001000";	-- 0x01D4
		when 000235 => D <= "1011000010111100";	-- 0x01D6
		when 000236 => D <= "0000000000000000";	-- 0x01D8
		when 000237 => D <= "0000000000000011";	-- 0x01DA
		when 000238 => D <= "0110011110100000";	-- 0x01DC
		when 000239 => D <= "0010011001111001";	-- 0x01DE
		when 000240 => D <= "0000000000000001";	-- 0x01E0
		when 000241 => D <= "0000000000100100";	-- 0x01E2
		when 000242 => D <= "0010110001001011";	-- 0x01E4
		when 000243 => D <= "1101011111000000";	-- 0x01E6
		when 000244 => D <= "0010000000111001";	-- 0x01E8
		when 000245 => D <= "0000000000000001";	-- 0x01EA
		when 000246 => D <= "0000000000101000";	-- 0x01EC
		when 000247 => D <= "1011000010001011";	-- 0x01EE
		when 000248 => D <= "0110001100000000";	-- 0x01F0
		when 000249 => D <= "0000100010000000";	-- 0x01F2
		when 000250 => D <= "0010001111001011";	-- 0x01F4
		when 000251 => D <= "0000000000000001";	-- 0x01F6
		when 000252 => D <= "0000000000100100";	-- 0x01F8
		when 000253 => D <= "0010001001001110";	-- 0x01FA
		when 000254 => D <= "0010010001001101";	-- 0x01FC
		when 000255 => D <= "0110000100000000";	-- 0x01FE
		when 000256 => D <= "0000100101110110";	-- 0x0200
		when 000257 => D <= "0010001001001000";	-- 0x0202
		when 000258 => D <= "0010010001001101";	-- 0x0204
		when 000259 => D <= "0010011001001100";	-- 0x0206
		when 000260 => D <= "0110000100000000";	-- 0x0208
		when 000261 => D <= "0000100101100000";	-- 0x020A
		when 000262 => D <= "0110000000000000";	-- 0x020C
		when 000263 => D <= "1111111101110000";	-- 0x020E
		when 000264 => D <= "0100110001001001";	-- 0x0210
		when 000265 => D <= "0101001111010100";	-- 0x0212
		when 000266 => D <= "0100110001001111";	-- 0x0214
		when 000267 => D <= "0100000111000100";	-- 0x0216
		when 000268 => D <= "0100111001000101";	-- 0x0218
		when 000269 => D <= "1101011101010010";	-- 0x021A
		when 000270 => D <= "0101010111001110";	-- 0x021C
		when 000271 => D <= "0101001101000001";	-- 0x021E
		when 000272 => D <= "0101011011000101";	-- 0x0220
		when 000273 => D <= "0100111001000101";	-- 0x0222
		when 000274 => D <= "0101100011010100";	-- 0x0224
		when 000275 => D <= "0100110001000101";	-- 0x0226
		when 000276 => D <= "1101010001001001";	-- 0x0228
		when 000277 => D <= "1100011001000111";	-- 0x022A
		when 000278 => D <= "0100111101010100";	-- 0x022C
		when 000279 => D <= "1100111101000111";	-- 0x022E
		when 000280 => D <= "0100111101010011";	-- 0x0230
		when 000281 => D <= "0101010111000010";	-- 0x0232
		when 000282 => D <= "0101001001000101";	-- 0x0234
		when 000283 => D <= "0101010001010101";	-- 0x0236
		when 000284 => D <= "0101001011001110";	-- 0x0238
		when 000285 => D <= "0101001001000101";	-- 0x023A
		when 000286 => D <= "1100110101000110";	-- 0x023C
		when 000287 => D <= "0100111111010010";	-- 0x023E
		when 000288 => D <= "0100100101001110";	-- 0x0240
		when 000289 => D <= "0101000001010101";	-- 0x0242
		when 000290 => D <= "1101010001010000";	-- 0x0244
		when 000291 => D <= "0101001001001001";	-- 0x0246
		when 000292 => D <= "0100111011010100";	-- 0x0248
		when 000293 => D <= "0101000001001111";	-- 0x024A
		when 000294 => D <= "0100101111000101";	-- 0x024C
		when 000295 => D <= "0101001101010100";	-- 0x024E
		when 000296 => D <= "0100111111010000";	-- 0x0250
		when 000297 => D <= "0100001001011001";	-- 0x0252
		when 000298 => D <= "1100010101000011";	-- 0x0254
		when 000299 => D <= "0100000101001100";	-- 0x0256
		when 000300 => D <= "1100110000000000";	-- 0x0258
		when 000301 => D <= "0101000001000101";	-- 0x025A
		when 000302 => D <= "0100010111001011";	-- 0x025C
		when 000303 => D <= "0101001001001110";	-- 0x025E
		when 000304 => D <= "1100010001000001";	-- 0x0260
		when 000305 => D <= "0100001011010011";	-- 0x0262
		when 000306 => D <= "0101001101001001";	-- 0x0264
		when 000307 => D <= "0101101011000101";	-- 0x0266
		when 000308 => D <= "0000000001010100";	-- 0x0268
		when 000309 => D <= "1100111100000000";	-- 0x026A
		when 000310 => D <= "0101001101010100";	-- 0x026C
		when 000311 => D <= "0100010111010000";	-- 0x026E
		when 000312 => D <= "0000000000111110";	-- 0x0270
		when 000313 => D <= "1011110100111100";	-- 0x0272
		when 000314 => D <= "1011111010111110";	-- 0x0274
		when 000315 => D <= "1011110100111100";	-- 0x0276
		when 000316 => D <= "1011110110111100";	-- 0x0278
		when 000317 => D <= "0000000000000000";	-- 0x027A
		when 000318 => D <= "0000000000000000";	-- 0x027C
		when 000319 => D <= "0000001111000000";	-- 0x027E
		when 000320 => D <= "0000000000000000";	-- 0x0280
		when 000321 => D <= "0000011001010010";	-- 0x0282
		when 000322 => D <= "0000000000000000";	-- 0x0284
		when 000323 => D <= "0000001101011010";	-- 0x0286
		when 000324 => D <= "0000000000000000";	-- 0x0288
		when 000325 => D <= "0000001101101110";	-- 0x028A
		when 000326 => D <= "0000000000000000";	-- 0x028C
		when 000327 => D <= "0000011010111010";	-- 0x028E
		when 000328 => D <= "0000000000000000";	-- 0x0290
		when 000329 => D <= "0000010100110100";	-- 0x0292
		when 000330 => D <= "0000000000000000";	-- 0x0294
		when 000331 => D <= "0000011001000010";	-- 0x0296
		when 000332 => D <= "0000000000000000";	-- 0x0298
		when 000333 => D <= "0000010110011010";	-- 0x029A
		when 000334 => D <= "0000000000000000";	-- 0x029C
		when 000335 => D <= "0000001110101100";	-- 0x029E
		when 000336 => D <= "0000000000000000";	-- 0x02A0
		when 000337 => D <= "0000010001100010";	-- 0x02A2
		when 000338 => D <= "0000000000000000";	-- 0x02A4
		when 000339 => D <= "0000010010010010";	-- 0x02A6
		when 000340 => D <= "0000000000000000";	-- 0x02A8
		when 000341 => D <= "0000010110010110";	-- 0x02AA
		when 000342 => D <= "0000000000000000";	-- 0x02AC
		when 000343 => D <= "0000010010110110";	-- 0x02AE
		when 000344 => D <= "0000000000000000";	-- 0x02B0
		when 000345 => D <= "0000010111000100";	-- 0x02B2
		when 000346 => D <= "0000000000000000";	-- 0x02B4
		when 000347 => D <= "0000001111110000";	-- 0x02B6
		when 000348 => D <= "0000000000000000";	-- 0x02B8
		when 000349 => D <= "0000011101000010";	-- 0x02BA
		when 000350 => D <= "0000000000000000";	-- 0x02BC
		when 000351 => D <= "0000001101100110";	-- 0x02BE
		when 000352 => D <= "0000000000000000";	-- 0x02C0
		when 000353 => D <= "0000000100011100";	-- 0x02C2
		when 000354 => D <= "0000000000000000";	-- 0x02C4
		when 000355 => D <= "0000011101011110";	-- 0x02C6
		when 000356 => D <= "0000000000000000";	-- 0x02C8
		when 000357 => D <= "0000011000111010";	-- 0x02CA
		when 000358 => D <= "0000000000000000";	-- 0x02CC
		when 000359 => D <= "0000100110000000";	-- 0x02CE
		when 000360 => D <= "0000000000000000";	-- 0x02D0
		when 000361 => D <= "0000100110001100";	-- 0x02D2
		when 000362 => D <= "0000000000000000";	-- 0x02D4
		when 000363 => D <= "0000100111000110";	-- 0x02D6
		when 000364 => D <= "0000000000000000";	-- 0x02D8
		when 000365 => D <= "0000100111011000";	-- 0x02DA
		when 000366 => D <= "0000000000000000";	-- 0x02DC
		when 000367 => D <= "0000100001101000";	-- 0x02DE
		when 000368 => D <= "0000000000000000";	-- 0x02E0
		when 000369 => D <= "0000010011010000";	-- 0x02E2
		when 000370 => D <= "0000000000000000";	-- 0x02E4
		when 000371 => D <= "0000101000101100";	-- 0x02E6
		when 000372 => D <= "0000000000000000";	-- 0x02E8
		when 000373 => D <= "0000010011100110";	-- 0x02EA
		when 000374 => D <= "0000000000000000";	-- 0x02EC
		when 000375 => D <= "0000010011101110";	-- 0x02EE
		when 000376 => D <= "0000000000000000";	-- 0x02F0
		when 000377 => D <= "0000011110000110";	-- 0x02F2
		when 000378 => D <= "0000000000000000";	-- 0x02F4
		when 000379 => D <= "0000011110010010";	-- 0x02F6
		when 000380 => D <= "0000000000000000";	-- 0x02F8
		when 000381 => D <= "0000011110011110";	-- 0x02FA
		when 000382 => D <= "0000000000000000";	-- 0x02FC
		when 000383 => D <= "0000011110110110";	-- 0x02FE
		when 000384 => D <= "0000000000000000";	-- 0x0300
		when 000385 => D <= "0000011110101010";	-- 0x0302
		when 000386 => D <= "0000000000000000";	-- 0x0304
		when 000387 => D <= "0000011111000100";	-- 0x0306
		when 000388 => D <= "0000000000000000";	-- 0x0308
		when 000389 => D <= "0000011111011010";	-- 0x030A
		when 000390 => D <= "0100001111111000";	-- 0x030C
		when 000391 => D <= "0000001000010000";	-- 0x030E
		when 000392 => D <= "0100010111111000";	-- 0x0310
		when 000393 => D <= "0000001001111100";	-- 0x0312
		when 000394 => D <= "0110000100000000";	-- 0x0314
		when 000395 => D <= "0000101000010010";	-- 0x0316
		when 000396 => D <= "0010011001001000";	-- 0x0318
		when 000397 => D <= "0100001000000010";	-- 0x031A
		when 000398 => D <= "0001000000011000";	-- 0x031C
		when 000399 => D <= "0001001000010001";	-- 0x031E
		when 000400 => D <= "0110011000000000";	-- 0x0320
		when 000401 => D <= "0000000000001000";	-- 0x0322
		when 000402 => D <= "0010000001001011";	-- 0x0324
		when 000403 => D <= "0110000000000000";	-- 0x0326
		when 000404 => D <= "0000000000101010";	-- 0x0328
		when 000405 => D <= "0001011000000000";	-- 0x032A
		when 000406 => D <= "1100011000000010";	-- 0x032C
		when 000407 => D <= "1011011000111100";	-- 0x032E
		when 000408 => D <= "0000000000101110";	-- 0x0330
		when 000409 => D <= "0110011100000000";	-- 0x0332
		when 000410 => D <= "0000000000011110";	-- 0x0334
		when 000411 => D <= "1100001000111100";	-- 0x0336
		when 000412 => D <= "0000000001111111";	-- 0x0338
		when 000413 => D <= "1011001000000000";	-- 0x033A
		when 000414 => D <= "0110011100000000";	-- 0x033C
		when 000415 => D <= "0000000000001110";	-- 0x033E
		when 000416 => D <= "0101100010001010";	-- 0x0340
		when 000417 => D <= "0010000001001011";	-- 0x0342
		when 000418 => D <= "0100001000000010";	-- 0x0344
		when 000419 => D <= "0100101000011001";	-- 0x0346
		when 000420 => D <= "0110101011111100";	-- 0x0348
		when 000421 => D <= "0110000011010000";	-- 0x034A
		when 000422 => D <= "0111010011111111";	-- 0x034C
		when 000423 => D <= "0100101000011001";	-- 0x034E
		when 000424 => D <= "0110101011001010";	-- 0x0350
		when 000425 => D <= "0100011111111000";	-- 0x0352
		when 000426 => D <= "0000000000000000";	-- 0x0354
		when 000427 => D <= "0010011001010010";	-- 0x0356
		when 000428 => D <= "0100111011010011";	-- 0x0358
		when 000429 => D <= "0110000100000000";	-- 0x035A
		when 000430 => D <= "0000011011000010";	-- 0x035C
		when 000431 => D <= "0010001111111000";	-- 0x035E
		when 000432 => D <= "0000000100000000";	-- 0x0360
		when 000433 => D <= "0000000000000001";	-- 0x0362
		when 000434 => D <= "0000000000100100";	-- 0x0364
		when 000435 => D <= "0110000100000000";	-- 0x0366
		when 000436 => D <= "0000011010110110";	-- 0x0368
		when 000437 => D <= "0110000000000000";	-- 0x036A
		when 000438 => D <= "1111110111110000";	-- 0x036C
		when 000439 => D <= "0110000100000000";	-- 0x036E
		when 000440 => D <= "0000011010101110";	-- 0x0370
		when 000441 => D <= "0010000001111000";	-- 0x0372
		when 000442 => D <= "0000000100000000";	-- 0x0374
		when 000443 => D <= "0010001111001000";	-- 0x0376
		when 000444 => D <= "0000000000000001";	-- 0x0378
		when 000445 => D <= "0000000000000100";	-- 0x037A
		when 000446 => D <= "0100101010111001";	-- 0x037C
		when 000447 => D <= "0000000000000001";	-- 0x037E
		when 000448 => D <= "0000000000000100";	-- 0x0380
		when 000449 => D <= "0110011100000000";	-- 0x0382
		when 000450 => D <= "1111110111011000";	-- 0x0384
		when 000451 => D <= "0100001010000001";	-- 0x0386
		when 000452 => D <= "0010001001001000";	-- 0x0388
		when 000453 => D <= "0110000100000000";	-- 0x038A
		when 000454 => D <= "0000011110110110";	-- 0x038C
		when 000455 => D <= "0110010100000000";	-- 0x038E
		when 000456 => D <= "1111110111001100";	-- 0x0390
		when 000457 => D <= "0010001111001001";	-- 0x0392
		when 000458 => D <= "0000000000000001";	-- 0x0394
		when 000459 => D <= "0000000000000100";	-- 0x0396
		when 000460 => D <= "0010000001001001";	-- 0x0398
		when 000461 => D <= "0101010010001000";	-- 0x039A
		when 000462 => D <= "0110000100000000";	-- 0x039C
		when 000463 => D <= "0000100111110010";	-- 0x039E
		when 000464 => D <= "0100001111111000";	-- 0x03A0
		when 000465 => D <= "0000001000100010";	-- 0x03A2
		when 000466 => D <= "0100010111111000";	-- 0x03A4
		when 000467 => D <= "0000001010010000";	-- 0x03A6
		when 000468 => D <= "0110000000000000";	-- 0x03A8
		when 000469 => D <= "1111111101101010";	-- 0x03AA
		when 000470 => D <= "0110000100000000";	-- 0x03AC
		when 000471 => D <= "0000001111000110";	-- 0x03AE
		when 000472 => D <= "0110000100000000";	-- 0x03B0
		when 000473 => D <= "0000011001101100";	-- 0x03B2
		when 000474 => D <= "0010001000000000";	-- 0x03B4
		when 000475 => D <= "0110000100000000";	-- 0x03B6
		when 000476 => D <= "0000011101111100";	-- 0x03B8
		when 000477 => D <= "0110011000000000";	-- 0x03BA
		when 000478 => D <= "0000011011000000";	-- 0x03BC
		when 000479 => D <= "0110000011010010";	-- 0x03BE
		when 000480 => D <= "0110000100000000";	-- 0x03C0
		when 000481 => D <= "0000100100101010";	-- 0x03C2
		when 000482 => D <= "0110000100000000";	-- 0x03C4
		when 000483 => D <= "0000011001011000";	-- 0x03C6
		when 000484 => D <= "0110000100000000";	-- 0x03C8
		when 000485 => D <= "0000011101101010";	-- 0x03CA
		when 000486 => D <= "0110010100000000";	-- 0x03CC
		when 000487 => D <= "1111110110001110";	-- 0x03CE
		when 000488 => D <= "0110000100000000";	-- 0x03D0
		when 000489 => D <= "0000100011100010";	-- 0x03D2
		when 000490 => D <= "0110000100000000";	-- 0x03D4
		when 000491 => D <= "0000100110111010";	-- 0x03D6
		when 000492 => D <= "0110011100000000";	-- 0x03D8
		when 000493 => D <= "0000000000010000";	-- 0x03DA
		when 000494 => D <= "1011000000111100";	-- 0x03DC
		when 000495 => D <= "0000000000010011";	-- 0x03DE
		when 000496 => D <= "0110011000000000";	-- 0x03E0
		when 000497 => D <= "0000000000001000";	-- 0x03E2
		when 000498 => D <= "0110000100000000";	-- 0x03E4
		when 000499 => D <= "0000100110101010";	-- 0x03E6
		when 000500 => D <= "0110011111111010";	-- 0x03E8
		when 000501 => D <= "0110000100000000";	-- 0x03EA
		when 000502 => D <= "0000011101010110";	-- 0x03EC
		when 000503 => D <= "0110000011011100";	-- 0x03EE
		when 000504 => D <= "0011100000111100";	-- 0x03F0
		when 000505 => D <= "0000000000001011";	-- 0x03F2
		when 000506 => D <= "0110000100000000";	-- 0x03F4
		when 000507 => D <= "0000100011011010";	-- 0x03F6
		when 000508 => D <= "0011101000000111";	-- 0x03F8
		when 000509 => D <= "0110000100000000";	-- 0x03FA
		when 000510 => D <= "0000100110101010";	-- 0x03FC
		when 000511 => D <= "0110000010011100";	-- 0x03FE
		when 000512 => D <= "0110000100000000";	-- 0x0400
		when 000513 => D <= "0000100011001110";	-- 0x0402
		when 000514 => D <= "0000110100001001";	-- 0x0404
		when 000515 => D <= "0110000100000000";	-- 0x0406
		when 000516 => D <= "0000100110011110";	-- 0x0408
		when 000517 => D <= "0110000000000000";	-- 0x040A
		when 000518 => D <= "1111111101110000";	-- 0x040C
		when 000519 => D <= "0110000100000000";	-- 0x040E
		when 000520 => D <= "0000100011000000";	-- 0x0410
		when 000521 => D <= "0010001100001011";	-- 0x0412
		when 000522 => D <= "0110000100000000";	-- 0x0414
		when 000523 => D <= "0000001101011110";	-- 0x0416
		when 000524 => D <= "0011100000000000";	-- 0x0418
		when 000525 => D <= "0110000000000000";	-- 0x041A
		when 000526 => D <= "0000000000011010";	-- 0x041C
		when 000527 => D <= "0110000100000000";	-- 0x041E
		when 000528 => D <= "0000100010110000";	-- 0x0420
		when 000529 => D <= "0010010000001101";	-- 0x0422
		when 000530 => D <= "0110000100000000";	-- 0x0424
		when 000531 => D <= "0000001101001110";	-- 0x0426
		when 000532 => D <= "0110000100000000";	-- 0x0428
		when 000533 => D <= "1111110011100010";	-- 0x042A
		when 000534 => D <= "0110000000000000";	-- 0x042C
		when 000535 => D <= "0000000000001000";	-- 0x042E
		when 000536 => D <= "0110000100000000";	-- 0x0430
		when 000537 => D <= "0000011111000100";	-- 0x0432
		when 000538 => D <= "0110000000010100";	-- 0x0434
		when 000539 => D <= "0110000100000000";	-- 0x0436
		when 000540 => D <= "0000100010011000";	-- 0x0438
		when 000541 => D <= "0010110000000111";	-- 0x043A
		when 000542 => D <= "0110000100000000";	-- 0x043C
		when 000543 => D <= "0000010111000110";	-- 0x043E
		when 000544 => D <= "0110000011001100";	-- 0x0440
		when 000545 => D <= "0110000100000000";	-- 0x0442
		when 000546 => D <= "0000100101100010";	-- 0x0444
		when 000547 => D <= "0110000000000000";	-- 0x0446
		when 000548 => D <= "0000000000010010";	-- 0x0448
		when 000549 => D <= "0011111100000100";	-- 0x044A
		when 000550 => D <= "0110000100000000";	-- 0x044C
		when 000551 => D <= "0000001100100110";	-- 0x044E
		when 000552 => D <= "0011100000011111";	-- 0x0450
		when 000553 => D <= "0010001000000000";	-- 0x0452
		when 000554 => D <= "0110000100000000";	-- 0x0454
		when 000555 => D <= "0000011111011110";	-- 0x0456
		when 000556 => D <= "0110000011011100";	-- 0x0458
		when 000557 => D <= "0110000100000000";	-- 0x045A
		when 000558 => D <= "0000010110101000";	-- 0x045C
		when 000559 => D <= "0110000000000000";	-- 0x045E
		when 000560 => D <= "0000010111001100";	-- 0x0460
		when 000561 => D <= "0110000100000000";	-- 0x0462
		when 000562 => D <= "0000011101000000";	-- 0x0464
		when 000563 => D <= "0110000100000000";	-- 0x0466
		when 000564 => D <= "0000001100001100";	-- 0x0468
		when 000565 => D <= "0010111100001000";	-- 0x046A
		when 000566 => D <= "0010001000000000";	-- 0x046C
		when 000567 => D <= "0110000100000000";	-- 0x046E
		when 000568 => D <= "0000011011000100";	-- 0x0470
		when 000569 => D <= "0110011000000000";	-- 0x0472
		when 000570 => D <= "0000011000001010";	-- 0x0474
		when 000571 => D <= "0010111100111001";	-- 0x0476
		when 000572 => D <= "0000000000000001";	-- 0x0478
		when 000573 => D <= "0000000000000100";	-- 0x047A
		when 000574 => D <= "0010111100111001";	-- 0x047C
		when 000575 => D <= "0000000000000001";	-- 0x047E
		when 000576 => D <= "0000000000001000";	-- 0x0480
		when 000577 => D <= "0100001010111001";	-- 0x0482
		when 000578 => D <= "0000000000000001";	-- 0x0484
		when 000579 => D <= "0000000000010000";	-- 0x0486
		when 000580 => D <= "0010001111001111";	-- 0x0488
		when 000581 => D <= "0000000000000001";	-- 0x048A
		when 000582 => D <= "0000000000001000";	-- 0x048C
		when 000583 => D <= "0110000000000000";	-- 0x048E
		when 000584 => D <= "1111111100000010";	-- 0x0490
		when 000585 => D <= "0110000100000000";	-- 0x0492
		when 000586 => D <= "0000010110001010";	-- 0x0494
		when 000587 => D <= "0010001000111001";	-- 0x0496
		when 000588 => D <= "0000000000000001";	-- 0x0498
		when 000589 => D <= "0000000000001000";	-- 0x049A
		when 000590 => D <= "0110011100000000";	-- 0x049C
		when 000591 => D <= "0000010110001110";	-- 0x049E
		when 000592 => D <= "0010111001000001";	-- 0x04A0
		when 000593 => D <= "0010001111011111";	-- 0x04A2
		when 000594 => D <= "0000000000000001";	-- 0x04A4
		when 000595 => D <= "0000000000001000";	-- 0x04A6
		when 000596 => D <= "0010001111011111";	-- 0x04A8
		when 000597 => D <= "0000000000000001";	-- 0x04AA
		when 000598 => D <= "0000000000000100";	-- 0x04AC
		when 000599 => D <= "0010000001011111";	-- 0x04AE
		when 000600 => D <= "0110000100000000";	-- 0x04B0
		when 000601 => D <= "0000011011001100";	-- 0x04B2
		when 000602 => D <= "0110000010100100";	-- 0x04B4
		when 000603 => D <= "0110000100000000";	-- 0x04B6
		when 000604 => D <= "0000011011101100";	-- 0x04B8
		when 000605 => D <= "0110000100000000";	-- 0x04BA
		when 000606 => D <= "0000010100101010";	-- 0x04BC
		when 000607 => D <= "0010001111001110";	-- 0x04BE
		when 000608 => D <= "0000000000000001";	-- 0x04C0
		when 000609 => D <= "0000000000010000";	-- 0x04C2
		when 000610 => D <= "0100001111111000";	-- 0x04C4
		when 000611 => D <= "0000001001101001";	-- 0x04C6
		when 000612 => D <= "0100010111111000";	-- 0x04C8
		when 000613 => D <= "0000001011100000";	-- 0x04CA
		when 000614 => D <= "0110000000000000";	-- 0x04CC
		when 000615 => D <= "1111111001000110";	-- 0x04CE
		when 000616 => D <= "0110000100000000";	-- 0x04D0
		when 000617 => D <= "0000001010100010";	-- 0x04D2
		when 000618 => D <= "0010001111000000";	-- 0x04D4
		when 000619 => D <= "0000000000000001";	-- 0x04D6
		when 000620 => D <= "0000000000011000";	-- 0x04D8
		when 000621 => D <= "0100001111111000";	-- 0x04DA
		when 000622 => D <= "0000001001101100";	-- 0x04DC
		when 000623 => D <= "0100010111111000";	-- 0x04DE
		when 000624 => D <= "0000001011101000";	-- 0x04E0
		when 000625 => D <= "0110000000000000";	-- 0x04E2
		when 000626 => D <= "1111111000110000";	-- 0x04E4
		when 000627 => D <= "0110000100000000";	-- 0x04E6
		when 000628 => D <= "0000001010001100";	-- 0x04E8
		when 000629 => D <= "0110000000000000";	-- 0x04EA
		when 000630 => D <= "0000000000000100";	-- 0x04EC
		when 000631 => D <= "0111000000000001";	-- 0x04EE
		when 000632 => D <= "0010001111000000";	-- 0x04F0
		when 000633 => D <= "0000000000000001";	-- 0x04F2
		when 000634 => D <= "0000000000010100";	-- 0x04F4
		when 000635 => D <= "0010001111111001";	-- 0x04F6
		when 000636 => D <= "0000000000000001";	-- 0x04F8
		when 000637 => D <= "0000000000000100";	-- 0x04FA
		when 000638 => D <= "0000000000000001";	-- 0x04FC
		when 000639 => D <= "0000000000011100";	-- 0x04FE
		when 000640 => D <= "0010001111001000";	-- 0x0500
		when 000641 => D <= "0000000000000001";	-- 0x0502
		when 000642 => D <= "0000000000100000";	-- 0x0504
		when 000643 => D <= "0010110001001111";	-- 0x0506
		when 000644 => D <= "0110000000000000";	-- 0x0508
		when 000645 => D <= "0000000000001000";	-- 0x050A
		when 000646 => D <= "1101110111111100";	-- 0x050C
		when 000647 => D <= "0000000000000000";	-- 0x050E
		when 000648 => D <= "0000000000010100";	-- 0x0510
		when 000649 => D <= "0010000000010110";	-- 0x0512
		when 000650 => D <= "0110011100000000";	-- 0x0514
		when 000651 => D <= "0000000000011010";	-- 0x0516
		when 000652 => D <= "1011000010111001";	-- 0x0518
		when 000653 => D <= "0000000000000001";	-- 0x051A
		when 000654 => D <= "0000000000010000";	-- 0x051C
		when 000655 => D <= "0110011011101100";	-- 0x051E
		when 000656 => D <= "0010010001001111";	-- 0x0520
		when 000657 => D <= "0010001001001110";	-- 0x0522
		when 000658 => D <= "0100011111111000";	-- 0x0524
		when 000659 => D <= "0000000000010100";	-- 0x0526
		when 000660 => D <= "1101011111001001";	-- 0x0528
		when 000661 => D <= "0110000100000000";	-- 0x052A
		when 000662 => D <= "0000011001001010";	-- 0x052C
		when 000663 => D <= "0010111001001011";	-- 0x052E
		when 000664 => D <= "0110000000000000";	-- 0x0530
		when 000665 => D <= "1111111100101000";	-- 0x0532
		when 000666 => D <= "0110000100000000";	-- 0x0534
		when 000667 => D <= "0000001101100010";	-- 0x0536
		when 000668 => D <= "0110010100000000";	-- 0x0538
		when 000669 => D <= "0000010011110010";	-- 0x053A
		when 000670 => D <= "0010001001000000";	-- 0x053C
		when 000671 => D <= "0010000000111001";	-- 0x053E
		when 000672 => D <= "0000000000000001";	-- 0x0540
		when 000673 => D <= "0000000000010000";	-- 0x0542
		when 000674 => D <= "0110011100000000";	-- 0x0544
		when 000675 => D <= "0000010011100110";	-- 0x0546
		when 000676 => D <= "1011001111000000";	-- 0x0548
		when 000677 => D <= "0110011100000000";	-- 0x054A
		when 000678 => D <= "0000000000001000";	-- 0x054C
		when 000679 => D <= "0110000100000000";	-- 0x054E
		when 000680 => D <= "0000011000101110";	-- 0x0550
		when 000681 => D <= "0110000011101010";	-- 0x0552
		when 000682 => D <= "0010000000010001";	-- 0x0554
		when 000683 => D <= "1101000010111001";	-- 0x0556
		when 000684 => D <= "0000000000000001";	-- 0x0558
		when 000685 => D <= "0000000000010100";	-- 0x055A
		when 000686 => D <= "0110100100000000";	-- 0x055C
		when 000687 => D <= "0000010100011110";	-- 0x055E
		when 000688 => D <= "0010001010000000";	-- 0x0560
		when 000689 => D <= "0010001000111001";	-- 0x0562
		when 000690 => D <= "0000000000000001";	-- 0x0564
		when 000691 => D <= "0000000000011000";	-- 0x0566
		when 000692 => D <= "0100101010111001";	-- 0x0568
		when 000693 => D <= "0000000000000001";	-- 0x056A
		when 000694 => D <= "0000000000010100";	-- 0x056C
		when 000695 => D <= "0110101000000000";	-- 0x056E
		when 000696 => D <= "0000000000000100";	-- 0x0570
		when 000697 => D <= "1100000101000001";	-- 0x0572
		when 000698 => D <= "1011001010000000";	-- 0x0574
		when 000699 => D <= "0110110100000000";	-- 0x0576
		when 000700 => D <= "0000000000010110";	-- 0x0578
		when 000701 => D <= "0010001111111001";	-- 0x057A
		when 000702 => D <= "0000000000000001";	-- 0x057C
		when 000703 => D <= "0000000000011100";	-- 0x057E
		when 000704 => D <= "0000000000000001";	-- 0x0580
		when 000705 => D <= "0000000000000100";	-- 0x0582
		when 000706 => D <= "0010000001111001";	-- 0x0584
		when 000707 => D <= "0000000000000001";	-- 0x0586
		when 000708 => D <= "0000000000100000";	-- 0x0588
		when 000709 => D <= "0110000000000000";	-- 0x058A
		when 000710 => D <= "1111111011001110";	-- 0x058C
		when 000711 => D <= "0110000100000000";	-- 0x058E
		when 000712 => D <= "0000010111101110";	-- 0x0590
		when 000713 => D <= "0110000000000000";	-- 0x0592
		when 000714 => D <= "1111111011000110";	-- 0x0594
		when 000715 => D <= "0110000000000000";	-- 0x0596
		when 000716 => D <= "0000000000001100";	-- 0x0598
		when 000717 => D <= "0110000100000000";	-- 0x059A
		when 000718 => D <= "0000000111011000";	-- 0x059C
		when 000719 => D <= "0100101010000000";	-- 0x059E
		when 000720 => D <= "0110011000000000";	-- 0x05A0
		when 000721 => D <= "1111110111111010";	-- 0x05A2
		when 000722 => D <= "0010001001001000";	-- 0x05A4
		when 000723 => D <= "0100001010000001";	-- 0x05A6
		when 000724 => D <= "0110000100000000";	-- 0x05A8
		when 000725 => D <= "0000010110111000";	-- 0x05AA
		when 000726 => D <= "0110010000000000";	-- 0x05AC
		when 000727 => D <= "1111110111100100";	-- 0x05AE
		when 000728 => D <= "0110000000000000";	-- 0x05B0
		when 000729 => D <= "1111101110101010";	-- 0x05B2
		when 000730 => D <= "0010111001111001";	-- 0x05B4
		when 000731 => D <= "0000000000000001";	-- 0x05B6
		when 000732 => D <= "0000000000001100";	-- 0x05B8
		when 000733 => D <= "0010001111011111";	-- 0x05BA
		when 000734 => D <= "0000000000000001";	-- 0x05BC
		when 000735 => D <= "0000000000000100";	-- 0x05BE
		when 000736 => D <= "0101100010001111";	-- 0x05C0
		when 000737 => D <= "0010000001011111";	-- 0x05C2
		when 000738 => D <= "0010111100001000";	-- 0x05C4
		when 000739 => D <= "0110000100000000";	-- 0x05C6
		when 000740 => D <= "0000011000101110";	-- 0x05C8
		when 000741 => D <= "0110000000001110";	-- 0x05CA
		when 000742 => D <= "0110000100000000";	-- 0x05CC
		when 000743 => D <= "0000001011001010";	-- 0x05CE
		when 000744 => D <= "0110010100000000";	-- 0x05D0
		when 000745 => D <= "0000000001011010";	-- 0x05D2
		when 000746 => D <= "0010010001000000";	-- 0x05D4
		when 000747 => D <= "0110000000000000";	-- 0x05D6
		when 000748 => D <= "0000000000011100";	-- 0x05D8
		when 000749 => D <= "0010111100001000";	-- 0x05DA
		when 000750 => D <= "0110000100000000";	-- 0x05DC
		when 000751 => D <= "0000001010111010";	-- 0x05DE
		when 000752 => D <= "0110010100000000";	-- 0x05E0
		when 000753 => D <= "0000010001001010";	-- 0x05E2
		when 000754 => D <= "0010010001000000";	-- 0x05E4
		when 000755 => D <= "0001010000010000";	-- 0x05E6
		when 000756 => D <= "0100001000000000";	-- 0x05E8
		when 000757 => D <= "0001000010000000";	-- 0x05EA
		when 000758 => D <= "0010001001011111";	-- 0x05EC
		when 000759 => D <= "0110000100000000";	-- 0x05EE
		when 000760 => D <= "0000010111101000";	-- 0x05F0
		when 000761 => D <= "0001000010000010";	-- 0x05F2
		when 000762 => D <= "0010111100001000";	-- 0x05F4
		when 000763 => D <= "0010111100111001";	-- 0x05F6
		when 000764 => D <= "0000000000000001";	-- 0x05F8
		when 000765 => D <= "0000000000000100";	-- 0x05FA
		when 000766 => D <= "0010001111111100";	-- 0x05FC
		when 000767 => D <= "1111111111111111";	-- 0x05FE
		when 000768 => D <= "1111111111111111";	-- 0x0600
		when 000769 => D <= "0000000000000001";	-- 0x0602
		when 000770 => D <= "0000000000000100";	-- 0x0604
		when 000771 => D <= "0010001111001111";	-- 0x0606
		when 000772 => D <= "0000000000000001";	-- 0x0608
		when 000773 => D <= "0000000000001100";	-- 0x060A
		when 000774 => D <= "0010111100001010";	-- 0x060C
		when 000775 => D <= "0001000000111100";	-- 0x060E
		when 000776 => D <= "0000000000111010";	-- 0x0610
		when 000777 => D <= "0110000100000000";	-- 0x0612
		when 000778 => D <= "0000010001110010";	-- 0x0614
		when 000779 => D <= "0100000111111001";	-- 0x0616
		when 000780 => D <= "0000000000000001";	-- 0x0618
		when 000781 => D <= "0000000000110000";	-- 0x061A
		when 000782 => D <= "0110000100000000";	-- 0x061C
		when 000783 => D <= "0000000101010110";	-- 0x061E
		when 000784 => D <= "0010010001011111";	-- 0x0620
		when 000785 => D <= "0010010010000000";	-- 0x0622
		when 000786 => D <= "0010001111011111";	-- 0x0624
		when 000787 => D <= "0000000000000001";	-- 0x0626
		when 000788 => D <= "0000000000000100";	-- 0x0628
		when 000789 => D <= "0010000001011111";	-- 0x062A
		when 000790 => D <= "0101100010001111";	-- 0x062C
		when 000791 => D <= "0110000100000000";	-- 0x062E
		when 000792 => D <= "0000011010100000";	-- 0x0630
		when 000793 => D <= "0010110000000011";	-- 0x0632
		when 000794 => D <= "0110000010001110";	-- 0x0634
		when 000795 => D <= "0110000000000000";	-- 0x0636
		when 000796 => D <= "1111111000100010";	-- 0x0638
		when 000797 => D <= "0000110000010000";	-- 0x063A
		when 000798 => D <= "0000000000001101";	-- 0x063C
		when 000799 => D <= "0110011100000000";	-- 0x063E
		when 000800 => D <= "0000000000001110";	-- 0x0640
		when 000801 => D <= "0110000100000000";	-- 0x0642
		when 000802 => D <= "0000001110100010";	-- 0x0644
		when 000803 => D <= "0110000100000000";	-- 0x0646
		when 000804 => D <= "0000011010001000";	-- 0x0648
		when 000805 => D <= "0010110000000011";	-- 0x064A
		when 000806 => D <= "0110000011110100";	-- 0x064C
		when 000807 => D <= "0110000000000000";	-- 0x064E
		when 000808 => D <= "1111111000001010";	-- 0x0650
		when 000809 => D <= "0010000001111000";	-- 0x0652
		when 000810 => D <= "0000000100000000";	-- 0x0654
		when 000811 => D <= "0001000000111100";	-- 0x0656
		when 000812 => D <= "0000000000001101";	-- 0x0658
		when 000813 => D <= "0110000100000000";	-- 0x065A
		when 000814 => D <= "1111101010111000";	-- 0x065C
		when 000815 => D <= "0110000100000000";	-- 0x065E
		when 000816 => D <= "1111101010111000";	-- 0x0660
		when 000817 => D <= "0110011111111010";	-- 0x0662
		when 000818 => D <= "1011000000111100";	-- 0x0664
		when 000819 => D <= "0000000001000000";	-- 0x0666
		when 000820 => D <= "0110011100000000";	-- 0x0668
		when 000821 => D <= "0000000000100100";	-- 0x066A
		when 000822 => D <= "1011000000111100";	-- 0x066C
		when 000823 => D <= "0000000000111010";	-- 0x066E
		when 000824 => D <= "0110011011101100";	-- 0x0670
		when 000825 => D <= "0110000100000000";	-- 0x0672
		when 000826 => D <= "0000000000100100";	-- 0x0674
		when 000827 => D <= "0001000011000001";	-- 0x0676
		when 000828 => D <= "0110000100000000";	-- 0x0678
		when 000829 => D <= "0000000000011110";	-- 0x067A
		when 000830 => D <= "0001000011000001";	-- 0x067C
		when 000831 => D <= "0110000100000000";	-- 0x067E
		when 000832 => D <= "1111101010011000";	-- 0x0680
		when 000833 => D <= "0110011111111010";	-- 0x0682
		when 000834 => D <= "0001000011000000";	-- 0x0684
		when 000835 => D <= "1011000000111100";	-- 0x0686
		when 000836 => D <= "0000000000001101";	-- 0x0688
		when 000837 => D <= "0110011011110010";	-- 0x068A
		when 000838 => D <= "0110000011010000";	-- 0x068C
		when 000839 => D <= "0010001111001000";	-- 0x068E
		when 000840 => D <= "0000000000000001";	-- 0x0690
		when 000841 => D <= "0000000000100100";	-- 0x0692
		when 000842 => D <= "0110000000000000";	-- 0x0694
		when 000843 => D <= "1111101011000110";	-- 0x0696
		when 000844 => D <= "0111010000000001";	-- 0x0698
		when 000845 => D <= "0100001001000001";	-- 0x069A
		when 000846 => D <= "0110000100000000";	-- 0x069C
		when 000847 => D <= "1111101001111010";	-- 0x069E
		when 000848 => D <= "0110011111111010";	-- 0x06A0
		when 000849 => D <= "1011000000111100";	-- 0x06A2
		when 000850 => D <= "0000000001000001";	-- 0x06A4
		when 000851 => D <= "0110010100000000";	-- 0x06A6
		when 000852 => D <= "0000000000000100";	-- 0x06A8
		when 000853 => D <= "0101111100000000";	-- 0x06AA
		when 000854 => D <= "1100000000111100";	-- 0x06AC
		when 000855 => D <= "0000000000001111";	-- 0x06AE
		when 000856 => D <= "1110100100001001";	-- 0x06B0
		when 000857 => D <= "1000001000000000";	-- 0x06B2
		when 000858 => D <= "0101000111001010";	-- 0x06B4
		when 000859 => D <= "1111111111100110";	-- 0x06B6
		when 000860 => D <= "0100111001110101";	-- 0x06B8
		when 000861 => D <= "0010000001111000";	-- 0x06BA
		when 000862 => D <= "0000000100000000";	-- 0x06BC
		when 000863 => D <= "0010001001111001";	-- 0x06BE
		when 000864 => D <= "0000000000000001";	-- 0x06C0
		when 000865 => D <= "0000000000100100";	-- 0x06C2
		when 000866 => D <= "0001000000111100";	-- 0x06C4
		when 000867 => D <= "0000000000001101";	-- 0x06C6
		when 000868 => D <= "0110000100000000";	-- 0x06C8
		when 000869 => D <= "1111101001001010";	-- 0x06CA
		when 000870 => D <= "0001000000111100";	-- 0x06CC
		when 000871 => D <= "0000000000001010";	-- 0x06CE
		when 000872 => D <= "0110000100000000";	-- 0x06D0
		when 000873 => D <= "1111101001000010";	-- 0x06D2
		when 000874 => D <= "1011001111001000";	-- 0x06D4
		when 000875 => D <= "0110001100000000";	-- 0x06D6
		when 000876 => D <= "0000000000100100";	-- 0x06D8
		when 000877 => D <= "0001000000111100";	-- 0x06DA
		when 000878 => D <= "0000000000111010";	-- 0x06DC
		when 000879 => D <= "0110000100000000";	-- 0x06DE
		when 000880 => D <= "1111101000110100";	-- 0x06E0
		when 000881 => D <= "0001001000011000";	-- 0x06E2
		when 000882 => D <= "0110000100000000";	-- 0x06E4
		when 000883 => D <= "0000000000111010";	-- 0x06E6
		when 000884 => D <= "0001001000011000";	-- 0x06E8
		when 000885 => D <= "0110000100000000";	-- 0x06EA
		when 000886 => D <= "0000000000110100";	-- 0x06EC
		when 000887 => D <= "0001000000011000";	-- 0x06EE
		when 000888 => D <= "1011000000111100";	-- 0x06F0
		when 000889 => D <= "0000000000001101";	-- 0x06F2
		when 000890 => D <= "0110011111001110";	-- 0x06F4
		when 000891 => D <= "0110000100000000";	-- 0x06F6
		when 000892 => D <= "1111101000011100";	-- 0x06F8
		when 000893 => D <= "0110000011110010";	-- 0x06FA
		when 000894 => D <= "0001000000111100";	-- 0x06FC
		when 000895 => D <= "0000000001000000";	-- 0x06FE
		when 000896 => D <= "0110000100000000";	-- 0x0700
		when 000897 => D <= "1111101000010010";	-- 0x0702
		when 000898 => D <= "0001000000111100";	-- 0x0704
		when 000899 => D <= "0000000000001101";	-- 0x0706
		when 000900 => D <= "0110000100000000";	-- 0x0708
		when 000901 => D <= "1111101000001010";	-- 0x070A
		when 000902 => D <= "0001000000111100";	-- 0x070C
		when 000903 => D <= "0000000000001010";	-- 0x070E
		when 000904 => D <= "0110000100000000";	-- 0x0710
		when 000905 => D <= "1111101000000010";	-- 0x0712
		when 000906 => D <= "0001000000111100";	-- 0x0714
		when 000907 => D <= "0000000000011010";	-- 0x0716
		when 000908 => D <= "0110000100000000";	-- 0x0718
		when 000909 => D <= "1111100111111010";	-- 0x071A
		when 000910 => D <= "0110000000000000";	-- 0x071C
		when 000911 => D <= "1111101000111110";	-- 0x071E
		when 000912 => D <= "0111010000000001";	-- 0x0720
		when 000913 => D <= "1110100100011001";	-- 0x0722
		when 000914 => D <= "0001000000000001";	-- 0x0724
		when 000915 => D <= "1100000000111100";	-- 0x0726
		when 000916 => D <= "0000000000001111";	-- 0x0728
		when 000917 => D <= "0000011000000000";	-- 0x072A
		when 000918 => D <= "0000000000110000";	-- 0x072C
		when 000919 => D <= "1011000000111100";	-- 0x072E
		when 000920 => D <= "0000000000111001";	-- 0x0730
		when 000921 => D <= "0110001100000000";	-- 0x0732
		when 000922 => D <= "0000000000000100";	-- 0x0734
		when 000923 => D <= "0101111000000000";	-- 0x0736
		when 000924 => D <= "0110000100000000";	-- 0x0738
		when 000925 => D <= "1111100111011010";	-- 0x073A
		when 000926 => D <= "0101000111001010";	-- 0x073C
		when 000927 => D <= "1111111111100100";	-- 0x073E
		when 000928 => D <= "0100111001110101";	-- 0x0740
		when 000929 => D <= "0110000100000000";	-- 0x0742
		when 000930 => D <= "0000000000110000";	-- 0x0744
		when 000931 => D <= "0110000100000000";	-- 0x0746
		when 000932 => D <= "0000010110001000";	-- 0x0748
		when 000933 => D <= "0010110000001111";	-- 0x074A
		when 000934 => D <= "0010111100000000";	-- 0x074C
		when 000935 => D <= "0110000100000000";	-- 0x074E
		when 000936 => D <= "0000000000100100";	-- 0x0750
		when 000937 => D <= "0010001001011111";	-- 0x0752
		when 000938 => D <= "0001001010000000";	-- 0x0754
		when 000939 => D <= "0110000000000000";	-- 0x0756
		when 000940 => D <= "1111110100000010";	-- 0x0758
		when 000941 => D <= "0110000000000000";	-- 0x075A
		when 000942 => D <= "0000001011010000";	-- 0x075C
		when 000943 => D <= "0110000100000000";	-- 0x075E
		when 000944 => D <= "0000000000010100";	-- 0x0760
		when 000945 => D <= "0100101010000000";	-- 0x0762
		when 000946 => D <= "0110011100000000";	-- 0x0764
		when 000947 => D <= "0000001100010110";	-- 0x0766
		when 000948 => D <= "0010111100001000";	-- 0x0768
		when 000949 => D <= "0010001001000000";	-- 0x076A
		when 000950 => D <= "0100111010010001";	-- 0x076C
		when 000951 => D <= "0010000001011111";	-- 0x076E
		when 000952 => D <= "0110000000000000";	-- 0x0770
		when 000953 => D <= "1111110011101000";	-- 0x0772
		when 000954 => D <= "0110000100000000";	-- 0x0774
		when 000955 => D <= "0000000001111010";	-- 0x0776
		when 000956 => D <= "0010111100000000";	-- 0x0778
		when 000957 => D <= "0100001111111000";	-- 0x077A
		when 000958 => D <= "0000001001110001";	-- 0x077C
		when 000959 => D <= "0100010111111000";	-- 0x077E
		when 000960 => D <= "0000001011110000";	-- 0x0780
		when 000961 => D <= "0110000000000000";	-- 0x0782
		when 000962 => D <= "1111101110010000";	-- 0x0784
		when 000963 => D <= "0110000100000000";	-- 0x0786
		when 000964 => D <= "0000000001010110";	-- 0x0788
		when 000965 => D <= "0110110100000000";	-- 0x078A
		when 000966 => D <= "0000000001000110";	-- 0x078C
		when 000967 => D <= "0110000000000000";	-- 0x078E
		when 000968 => D <= "0000000001000110";	-- 0x0790
		when 000969 => D <= "0110000100000000";	-- 0x0792
		when 000970 => D <= "0000000001001010";	-- 0x0794
		when 000971 => D <= "0110011100000000";	-- 0x0796
		when 000972 => D <= "0000000000111010";	-- 0x0798
		when 000973 => D <= "0110000000000000";	-- 0x079A
		when 000974 => D <= "0000000000111010";	-- 0x079C
		when 000975 => D <= "0110000100000000";	-- 0x079E
		when 000976 => D <= "0000000000111110";	-- 0x07A0
		when 000977 => D <= "0110111100000000";	-- 0x07A2
		when 000978 => D <= "0000000000101110";	-- 0x07A4
		when 000979 => D <= "0110000000000000";	-- 0x07A6
		when 000980 => D <= "0000000000101110";	-- 0x07A8
		when 000981 => D <= "0110000100000000";	-- 0x07AA
		when 000982 => D <= "0000000000110010";	-- 0x07AC
		when 000983 => D <= "0110111000000000";	-- 0x07AE
		when 000984 => D <= "0000000000100010";	-- 0x07B0
		when 000985 => D <= "0110000000000000";	-- 0x07B2
		when 000986 => D <= "0000000000100010";	-- 0x07B4
		when 000987 => D <= "0110000100000000";	-- 0x07B6
		when 000988 => D <= "0000000000100110";	-- 0x07B8
		when 000989 => D <= "0110011000000000";	-- 0x07BA
		when 000990 => D <= "0000000000010110";	-- 0x07BC
		when 000991 => D <= "0110000000000000";	-- 0x07BE
		when 000992 => D <= "0000000000010110";	-- 0x07C0
		when 000993 => D <= "0100111001110101";	-- 0x07C2
		when 000994 => D <= "0110000100000000";	-- 0x07C4
		when 000995 => D <= "0000000000011000";	-- 0x07C6
		when 000996 => D <= "0110110000000000";	-- 0x07C8
		when 000997 => D <= "0000000000001000";	-- 0x07CA
		when 000998 => D <= "0110000000000000";	-- 0x07CC
		when 000999 => D <= "0000000000001000";	-- 0x07CE
		when 001000 => D <= "0100111001110101";	-- 0x07D0
		when 001001 => D <= "0100001010000000";	-- 0x07D2
		when 001002 => D <= "0100111001110101";	-- 0x07D4
		when 001003 => D <= "0111000000000001";	-- 0x07D6
		when 001004 => D <= "0100111001110101";	-- 0x07D8
		when 001005 => D <= "0010000000011111";	-- 0x07DA
		when 001006 => D <= "0100111001110101";	-- 0x07DC
		when 001007 => D <= "0010000000011111";	-- 0x07DE
		when 001008 => D <= "0010001000011111";	-- 0x07E0
		when 001009 => D <= "0010111100000000";	-- 0x07E2
		when 001010 => D <= "0010111100000001";	-- 0x07E4
		when 001011 => D <= "0110000100000000";	-- 0x07E6
		when 001012 => D <= "0000000000001000";	-- 0x07E8
		when 001013 => D <= "0010001000011111";	-- 0x07EA
		when 001014 => D <= "1011001010000000";	-- 0x07EC
		when 001015 => D <= "0100111001110101";	-- 0x07EE
		when 001016 => D <= "0110000100000000";	-- 0x07F0
		when 001017 => D <= "0000010011011110";	-- 0x07F2
		when 001018 => D <= "0010110100000111";	-- 0x07F4
		when 001019 => D <= "0100001010000000";	-- 0x07F6
		when 001020 => D <= "0110000000000000";	-- 0x07F8
		when 001021 => D <= "0000000000101000";	-- 0x07FA
		when 001022 => D <= "0110000100000000";	-- 0x07FC
		when 001023 => D <= "0000010011010010";	-- 0x07FE
		when 001024 => D <= "0010101100000001";	-- 0x0800
		when 001025 => D <= "0110000100000000";	-- 0x0802
		when 001026 => D <= "0000000000101010";	-- 0x0804
		when 001027 => D <= "0110000100000000";	-- 0x0806
		when 001028 => D <= "0000010011001000";	-- 0x0808
		when 001029 => D <= "0010101100010001";	-- 0x080A
		when 001030 => D <= "0010111100000000";	-- 0x080C
		when 001031 => D <= "0110000100000000";	-- 0x080E
		when 001032 => D <= "0000000000011110";	-- 0x0810
		when 001033 => D <= "0010001000011111";	-- 0x0812
		when 001034 => D <= "1101000010000001";	-- 0x0814
		when 001035 => D <= "0110100100000000";	-- 0x0816
		when 001036 => D <= "0000001001100100";	-- 0x0818
		when 001037 => D <= "0110000011101010";	-- 0x081A
		when 001038 => D <= "0110000100000000";	-- 0x081C
		when 001039 => D <= "0000010010110010";	-- 0x081E
		when 001040 => D <= "0010110101110001";	-- 0x0820
		when 001041 => D <= "0010111100000000";	-- 0x0822
		when 001042 => D <= "0110000100000000";	-- 0x0824
		when 001043 => D <= "0000000000001000";	-- 0x0826
		when 001044 => D <= "0100010010000000";	-- 0x0828
		when 001045 => D <= "0100111011111000";	-- 0x082A
		when 001046 => D <= "0000100000010010";	-- 0x082C
		when 001047 => D <= "0110000100000000";	-- 0x082E
		when 001048 => D <= "0000000000101100";	-- 0x0830
		when 001049 => D <= "0110000100000000";	-- 0x0832
		when 001050 => D <= "0000010010011100";	-- 0x0834
		when 001051 => D <= "0010101000001111";	-- 0x0836
		when 001052 => D <= "0010111100000000";	-- 0x0838
		when 001053 => D <= "0110000100000000";	-- 0x083A
		when 001054 => D <= "0000000000100000";	-- 0x083C
		when 001055 => D <= "0010001000011111";	-- 0x083E
		when 001056 => D <= "0110000100000000";	-- 0x0840
		when 001057 => D <= "0000000010101110";	-- 0x0842
		when 001058 => D <= "0110000011101100";	-- 0x0844
		when 001059 => D <= "0110000100000000";	-- 0x0846
		when 001060 => D <= "0000010010001000";	-- 0x0848
		when 001061 => D <= "0010111101000111";	-- 0x084A
		when 001062 => D <= "0010111100000000";	-- 0x084C
		when 001063 => D <= "0110000100000000";	-- 0x084E
		when 001064 => D <= "0000000000001100";	-- 0x0850
		when 001065 => D <= "0010001000011111";	-- 0x0852
		when 001066 => D <= "1100000101000001";	-- 0x0854
		when 001067 => D <= "0110000100000000";	-- 0x0856
		when 001068 => D <= "0000000011100010";	-- 0x0858
		when 001069 => D <= "0110000011010110";	-- 0x085A
		when 001070 => D <= "0100001111111000";	-- 0x085C
		when 001071 => D <= "0000001001011010";	-- 0x085E
		when 001072 => D <= "0100010111111000";	-- 0x0860
		when 001073 => D <= "0000001011001100";	-- 0x0862
		when 001074 => D <= "0110000000000000";	-- 0x0864
		when 001075 => D <= "1111101010101110";	-- 0x0866
		when 001076 => D <= "0110000100000000";	-- 0x0868
		when 001077 => D <= "0000000000101110";	-- 0x086A
		when 001078 => D <= "0110010100000000";	-- 0x086C
		when 001079 => D <= "0000000000001010";	-- 0x086E
		when 001080 => D <= "0010001001000000";	-- 0x0870
		when 001081 => D <= "0100001010000000";	-- 0x0872
		when 001082 => D <= "0010000000010001";	-- 0x0874
		when 001083 => D <= "0100111001110101";	-- 0x0876
		when 001084 => D <= "0110000100000000";	-- 0x0878
		when 001085 => D <= "0000010001110010";	-- 0x087A
		when 001086 => D <= "0010000000000001";	-- 0x087C
		when 001087 => D <= "0100101001000010";	-- 0x087E
		when 001088 => D <= "0110011011110100";	-- 0x0880
		when 001089 => D <= "0110000100000000";	-- 0x0882
		when 001090 => D <= "0000010001001100";	-- 0x0884
		when 001091 => D <= "0010100000001101";	-- 0x0886
		when 001092 => D <= "0110000100000000";	-- 0x0888
		when 001093 => D <= "1111111011101010";	-- 0x088A
		when 001094 => D <= "0110000100000000";	-- 0x088C
		when 001095 => D <= "0000010001000010";	-- 0x088E
		when 001096 => D <= "0010100100000011";	-- 0x0890
		when 001097 => D <= "0100111001110101";	-- 0x0892
		when 001098 => D <= "0110000000000000";	-- 0x0894
		when 001099 => D <= "0000000110010110";	-- 0x0896
		when 001100 => D <= "0110000100000000";	-- 0x0898
		when 001101 => D <= "0000010010001110";	-- 0x089A
		when 001102 => D <= "0100001010000000";	-- 0x089C
		when 001103 => D <= "0001000000010000";	-- 0x089E
		when 001104 => D <= "0000010000000000";	-- 0x08A0
		when 001105 => D <= "0000000001000000";	-- 0x08A2
		when 001106 => D <= "0110010100000000";	-- 0x08A4
		when 001107 => D <= "0000000001001000";	-- 0x08A6
		when 001108 => D <= "0110011000000000";	-- 0x08A8
		when 001109 => D <= "0000000000101010";	-- 0x08AA
		when 001110 => D <= "0101001001001000";	-- 0x08AC
		when 001111 => D <= "0110000111010010";	-- 0x08AE
		when 001112 => D <= "1101000010000000";	-- 0x08B0
		when 001113 => D <= "0110010100000000";	-- 0x08B2
		when 001114 => D <= "0000000111001000";	-- 0x08B4
		when 001115 => D <= "1101000010000000";	-- 0x08B6
		when 001116 => D <= "0110010100000000";	-- 0x08B8
		when 001117 => D <= "0000000111000010";	-- 0x08BA
		when 001118 => D <= "0010111100000000";	-- 0x08BC
		when 001119 => D <= "0110000100000000";	-- 0x08BE
		when 001120 => D <= "0000000100011000";	-- 0x08C0
		when 001121 => D <= "0010001000011111";	-- 0x08C2
		when 001122 => D <= "1011000010000001";	-- 0x08C4
		when 001123 => D <= "0110001100000000";	-- 0x08C6
		when 001124 => D <= "0000000110101010";	-- 0x08C8
		when 001125 => D <= "0010000000111001";	-- 0x08CA
		when 001126 => D <= "0000000000000001";	-- 0x08CC
		when 001127 => D <= "0000000000101000";	-- 0x08CE
		when 001128 => D <= "1001000010000001";	-- 0x08D0
		when 001129 => D <= "0100111001110101";	-- 0x08D2
		when 001130 => D <= "1011000000111100";	-- 0x08D4
		when 001131 => D <= "0000000000011011";	-- 0x08D6
		when 001132 => D <= "0000101000111100";	-- 0x08D8
		when 001133 => D <= "0000000000000001";	-- 0x08DA
		when 001134 => D <= "0110010100000000";	-- 0x08DC
		when 001135 => D <= "0000000000010000";	-- 0x08DE
		when 001136 => D <= "0101001001001000";	-- 0x08E0
		when 001137 => D <= "1101000001000000";	-- 0x08E2
		when 001138 => D <= "1101000001000000";	-- 0x08E4
		when 001139 => D <= "0010001000111001";	-- 0x08E6
		when 001140 => D <= "0000000000000001";	-- 0x08E8
		when 001141 => D <= "0000000000101000";	-- 0x08EA
		when 001142 => D <= "1101000010000001";	-- 0x08EC
		when 001143 => D <= "0100111001110101";	-- 0x08EE
		when 001144 => D <= "0010100000000001";	-- 0x08F0
		when 001145 => D <= "1011000110000100";	-- 0x08F2
		when 001146 => D <= "0100101010000000";	-- 0x08F4
		when 001147 => D <= "0110101000000000";	-- 0x08F6
		when 001148 => D <= "0000000000000100";	-- 0x08F8
		when 001149 => D <= "0100010010000000";	-- 0x08FA
		when 001150 => D <= "0100101010000001";	-- 0x08FC
		when 001151 => D <= "0110101000000000";	-- 0x08FE
		when 001152 => D <= "0000000000000100";	-- 0x0900
		when 001153 => D <= "0100010010000001";	-- 0x0902
		when 001154 => D <= "1011001010111100";	-- 0x0904
		when 001155 => D <= "0000000000000000";	-- 0x0906
		when 001156 => D <= "1111111111111111";	-- 0x0908
		when 001157 => D <= "0110001100000000";	-- 0x090A
		when 001158 => D <= "0000000000001110";	-- 0x090C
		when 001159 => D <= "1100000101000001";	-- 0x090E
		when 001160 => D <= "1011001010111100";	-- 0x0910
		when 001161 => D <= "0000000000000000";	-- 0x0912
		when 001162 => D <= "1111111111111111";	-- 0x0914
		when 001163 => D <= "0110001000000000";	-- 0x0916
		when 001164 => D <= "0000000101100100";	-- 0x0918
		when 001165 => D <= "0011010000000000";	-- 0x091A
		when 001166 => D <= "1100010011000001";	-- 0x091C
		when 001167 => D <= "0100100001000000";	-- 0x091E
		when 001168 => D <= "1100000011000001";	-- 0x0920
		when 001169 => D <= "0100100001000000";	-- 0x0922
		when 001170 => D <= "0100101001000000";	-- 0x0924
		when 001171 => D <= "0110011000000000";	-- 0x0926
		when 001172 => D <= "0000000101010100";	-- 0x0928
		when 001173 => D <= "1101000010000010";	-- 0x092A
		when 001174 => D <= "0110101100000000";	-- 0x092C
		when 001175 => D <= "0000000101001110";	-- 0x092E
		when 001176 => D <= "0100101010000100";	-- 0x0930
		when 001177 => D <= "0110101000000000";	-- 0x0932
		when 001178 => D <= "0000000000000100";	-- 0x0934
		when 001179 => D <= "0100010010000000";	-- 0x0936
		when 001180 => D <= "0100111001110101";	-- 0x0938
		when 001181 => D <= "0100101010000001";	-- 0x093A
		when 001182 => D <= "0110011100000000";	-- 0x093C
		when 001183 => D <= "0000000100111110";	-- 0x093E
		when 001184 => D <= "0010010000000001";	-- 0x0940
		when 001185 => D <= "0010100000000001";	-- 0x0942
		when 001186 => D <= "1011000110000100";	-- 0x0944
		when 001187 => D <= "0100101010000000";	-- 0x0946
		when 001188 => D <= "0110101000000000";	-- 0x0948
		when 001189 => D <= "0000000000000100";	-- 0x094A
		when 001190 => D <= "0100010010000000";	-- 0x094C
		when 001191 => D <= "0100101010000001";	-- 0x094E
		when 001192 => D <= "0110101000000000";	-- 0x0950
		when 001193 => D <= "0000000000000100";	-- 0x0952
		when 001194 => D <= "0100010010000001";	-- 0x0954
		when 001195 => D <= "0111011000011111";	-- 0x0956
		when 001196 => D <= "0010001000000000";	-- 0x0958
		when 001197 => D <= "0100001010000000";	-- 0x095A
		when 001198 => D <= "1101001010000001";	-- 0x095C
		when 001199 => D <= "1101000110000000";	-- 0x095E
		when 001200 => D <= "0110011100000000";	-- 0x0960
		when 001201 => D <= "0000000000001100";	-- 0x0962
		when 001202 => D <= "1011000010000010";	-- 0x0964
		when 001203 => D <= "0110101100000000";	-- 0x0966
		when 001204 => D <= "0000000000000110";	-- 0x0968
		when 001205 => D <= "0101001010000001";	-- 0x096A
		when 001206 => D <= "1001000010000010";	-- 0x096C
		when 001207 => D <= "0101000111001011";	-- 0x096E
		when 001208 => D <= "1111111111101100";	-- 0x0970
		when 001209 => D <= "1100000101000001";	-- 0x0972
		when 001210 => D <= "0100101010000100";	-- 0x0974
		when 001211 => D <= "0110101000000000";	-- 0x0976
		when 001212 => D <= "0000000000000110";	-- 0x0978
		when 001213 => D <= "0100010010000000";	-- 0x097A
		when 001214 => D <= "0100010010000001";	-- 0x097C
		when 001215 => D <= "0100111001110101";	-- 0x097E
		when 001216 => D <= "0110000100000000";	-- 0x0980
		when 001217 => D <= "1111111100000000";	-- 0x0982
		when 001218 => D <= "0010001001000000";	-- 0x0984
		when 001219 => D <= "0100001010000000";	-- 0x0986
		when 001220 => D <= "0001000000010001";	-- 0x0988
		when 001221 => D <= "0100111001110101";	-- 0x098A
		when 001222 => D <= "0110000100000000";	-- 0x098C
		when 001223 => D <= "1111111011110100";	-- 0x098E
		when 001224 => D <= "0100101010000000";	-- 0x0990
		when 001225 => D <= "0110011100000000";	-- 0x0992
		when 001226 => D <= "0000000011101000";	-- 0x0994
		when 001227 => D <= "0110101100000000";	-- 0x0996
		when 001228 => D <= "0000000011100100";	-- 0x0998
		when 001229 => D <= "0010001000000000";	-- 0x099A
		when 001230 => D <= "0010001001111001";	-- 0x099C
		when 001231 => D <= "0000000000000001";	-- 0x099E
		when 001232 => D <= "0000000000000000";	-- 0x09A0
		when 001233 => D <= "1011001111111100";	-- 0x09A2
		when 001234 => D <= "0000000000000000";	-- 0x09A4
		when 001235 => D <= "0000111001011010";	-- 0x09A6
		when 001236 => D <= "0110010100000000";	-- 0x09A8
		when 001237 => D <= "0000000000000110";	-- 0x09AA
		when 001238 => D <= "0100001111111000";	-- 0x09AC
		when 001239 => D <= "0000000100000100";	-- 0x09AE
		when 001240 => D <= "0010000000011001";	-- 0x09B0
		when 001241 => D <= "0000100010000000";	-- 0x09B2
		when 001242 => D <= "0000000000011111";	-- 0x09B4
		when 001243 => D <= "0010001111001001";	-- 0x09B6
		when 001244 => D <= "0000000000000001";	-- 0x09B8
		when 001245 => D <= "0000000000000000";	-- 0x09BA
		when 001246 => D <= "0110000100000000";	-- 0x09BC
		when 001247 => D <= "1111111101111100";	-- 0x09BE
		when 001248 => D <= "0010000000000001";	-- 0x09C0
		when 001249 => D <= "0101001010000000";	-- 0x09C2
		when 001250 => D <= "0100111001110101";	-- 0x09C4
		when 001251 => D <= "0110000100000000";	-- 0x09C6
		when 001252 => D <= "1111111010111010";	-- 0x09C8
		when 001253 => D <= "0100101010000000";	-- 0x09CA
		when 001254 => D <= "0110101000000000";	-- 0x09CC
		when 001255 => D <= "0000000000001000";	-- 0x09CE
		when 001256 => D <= "0100010010000000";	-- 0x09D0
		when 001257 => D <= "0110101100000000";	-- 0x09D2
		when 001258 => D <= "0000000010101000";	-- 0x09D4
		when 001259 => D <= "0100111001110101";	-- 0x09D6
		when 001260 => D <= "0010000000111001";	-- 0x09D8
		when 001261 => D <= "0000000000000001";	-- 0x09DA
		when 001262 => D <= "0000000000101000";	-- 0x09DC
		when 001263 => D <= "1001000010111001";	-- 0x09DE
		when 001264 => D <= "0000000000000001";	-- 0x09E0
		when 001265 => D <= "0000000000100100";	-- 0x09E2
		when 001266 => D <= "0100111001110101";	-- 0x09E4
		when 001267 => D <= "0110000100000000";	-- 0x09E6
		when 001268 => D <= "1111111010110000";	-- 0x09E8
		when 001269 => D <= "0110010100000000";	-- 0x09EA
		when 001270 => D <= "0000000001000000";	-- 0x09EC
		when 001271 => D <= "0010111100000000";	-- 0x09EE
		when 001272 => D <= "0110000100000000";	-- 0x09F0
		when 001273 => D <= "0000001011011110";	-- 0x09F2
		when 001274 => D <= "0011110100001011";	-- 0x09F4
		when 001275 => D <= "0110000100000000";	-- 0x09F6
		when 001276 => D <= "1111110101111100";	-- 0x09F8
		when 001277 => D <= "0010110001011111";	-- 0x09FA
		when 001278 => D <= "0010110010000000";	-- 0x09FC
		when 001279 => D <= "0100111001110101";	-- 0x09FE
		when 001280 => D <= "0110000000000000";	-- 0x0A00
		when 001281 => D <= "0000000000101010";	-- 0x0A02
		when 001282 => D <= "0110000100000000";	-- 0x0A04
		when 001283 => D <= "0000001011001010";	-- 0x0A06
		when 001284 => D <= "0011101000000111";	-- 0x0A08
		when 001285 => D <= "0101100010001111";	-- 0x0A0A
		when 001286 => D <= "0110000000000000";	-- 0x0A0C
		when 001287 => D <= "1111100110001110";	-- 0x0A0E
		when 001288 => D <= "0110000100000000";	-- 0x0A10
		when 001289 => D <= "0000001010111110";	-- 0x0A12
		when 001290 => D <= "0000110100000111";	-- 0x0A14
		when 001291 => D <= "0101100010001111";	-- 0x0A16
		when 001292 => D <= "0110000000000000";	-- 0x0A18
		when 001293 => D <= "1111100101100010";	-- 0x0A1A
		when 001294 => D <= "0100111001110101";	-- 0x0A1C
		when 001295 => D <= "0110000100000000";	-- 0x0A1E
		when 001296 => D <= "0000001100001000";	-- 0x0A20
		when 001297 => D <= "0000110000010000";	-- 0x0A22
		when 001298 => D <= "0000000000001101";	-- 0x0A24
		when 001299 => D <= "0110011000000000";	-- 0x0A26
		when 001300 => D <= "0000000000000100";	-- 0x0A28
		when 001301 => D <= "0100111001110101";	-- 0x0A2A
		when 001302 => D <= "0010111100001000";	-- 0x0A2C
		when 001303 => D <= "0100110111111001";	-- 0x0A2E
		when 001304 => D <= "0000000000000000";	-- 0x0A30
		when 001305 => D <= "0000111001001000";	-- 0x0A32
		when 001306 => D <= "0110000100000000";	-- 0x0A34
		when 001307 => D <= "0000001101110110";	-- 0x0A36
		when 001308 => D <= "0010000001011111";	-- 0x0A38
		when 001309 => D <= "0010000000111001";	-- 0x0A3A
		when 001310 => D <= "0000000000000001";	-- 0x0A3C
		when 001311 => D <= "0000000000000100";	-- 0x0A3E
		when 001312 => D <= "0110011100000000";	-- 0x0A40
		when 001313 => D <= "1111011100011010";	-- 0x0A42
		when 001314 => D <= "1011000010111100";	-- 0x0A44
		when 001315 => D <= "1111111111111111";	-- 0x0A46
		when 001316 => D <= "1111111111111111";	-- 0x0A48
		when 001317 => D <= "0110011100000000";	-- 0x0A4A
		when 001318 => D <= "1111101101101000";	-- 0x0A4C
		when 001319 => D <= "0001111100010000";	-- 0x0A4E
		when 001320 => D <= "0100001000010000";	-- 0x0A50
		when 001321 => D <= "0010001001111001";	-- 0x0A52
		when 001322 => D <= "0000000000000001";	-- 0x0A54
		when 001323 => D <= "0000000000000100";	-- 0x0A56
		when 001324 => D <= "0110000100000000";	-- 0x0A58
		when 001325 => D <= "0000001001011010";	-- 0x0A5A
		when 001326 => D <= "0001000010011111";	-- 0x0A5C
		when 001327 => D <= "0001000000111100";	-- 0x0A5E
		when 001328 => D <= "0000000000111111";	-- 0x0A60
		when 001329 => D <= "0110000100000000";	-- 0x0A62
		when 001330 => D <= "1111011010101000";	-- 0x0A64
		when 001331 => D <= "0100001001000000";	-- 0x0A66
		when 001332 => D <= "0101001110001001";	-- 0x0A68
		when 001333 => D <= "0110000100000000";	-- 0x0A6A
		when 001334 => D <= "0000000101101100";	-- 0x0A6C
		when 001335 => D <= "0110000000000000";	-- 0x0A6E
		when 001336 => D <= "1111011011101100";	-- 0x0A70
		when 001337 => D <= "0010111100001000";	-- 0x0A72
		when 001338 => D <= "0100110111111001";	-- 0x0A74
		when 001339 => D <= "0000000000000000";	-- 0x0A76
		when 001340 => D <= "0000111001010000";	-- 0x0A78
		when 001341 => D <= "0110000010111000";	-- 0x0A7A
		when 001342 => D <= "0010111100001000";	-- 0x0A7C
		when 001343 => D <= "0100110111111001";	-- 0x0A7E
		when 001344 => D <= "0000000000000000";	-- 0x0A80
		when 001345 => D <= "0000111001000001";	-- 0x0A82
		when 001346 => D <= "0110000010101110";	-- 0x0A84
		when 001347 => D <= "0110000100000000";	-- 0x0A86
		when 001348 => D <= "1111011010000100";	-- 0x0A88
		when 001349 => D <= "0001000000111100";	-- 0x0A8A
		when 001350 => D <= "0000000000100000";	-- 0x0A8C
		when 001351 => D <= "0110000100000000";	-- 0x0A8E
		when 001352 => D <= "1111011001111100";	-- 0x0A90
		when 001353 => D <= "0100000111111001";	-- 0x0A92
		when 001354 => D <= "0000000000000001";	-- 0x0A94
		when 001355 => D <= "0000000000110000";	-- 0x0A96
		when 001356 => D <= "0110000100000000";	-- 0x0A98
		when 001357 => D <= "0000001011110110";	-- 0x0A9A
		when 001358 => D <= "0110011111111010";	-- 0x0A9C
		when 001359 => D <= "1011000000111100";	-- 0x0A9E
		when 001360 => D <= "0000000000001000";	-- 0x0AA0
		when 001361 => D <= "0110011100000000";	-- 0x0AA2
		when 001362 => D <= "0000000000101110";	-- 0x0AA4
		when 001363 => D <= "1011000000111100";	-- 0x0AA6
		when 001364 => D <= "0000000000011000";	-- 0x0AA8
		when 001365 => D <= "0110011100000000";	-- 0x0AAA
		when 001366 => D <= "0000000001001010";	-- 0x0AAC
		when 001367 => D <= "1011000000111100";	-- 0x0AAE
		when 001368 => D <= "0000000000001101";	-- 0x0AB0
		when 001369 => D <= "0110011100000000";	-- 0x0AB2
		when 001370 => D <= "0000000000001000";	-- 0x0AB4
		when 001371 => D <= "1011000000111100";	-- 0x0AB6
		when 001372 => D <= "0000000000100000";	-- 0x0AB8
		when 001373 => D <= "0110010111011100";	-- 0x0ABA
		when 001374 => D <= "0001000011000000";	-- 0x0ABC
		when 001375 => D <= "0110000100000000";	-- 0x0ABE
		when 001376 => D <= "1111011001001100";	-- 0x0AC0
		when 001377 => D <= "1011000000111100";	-- 0x0AC2
		when 001378 => D <= "0000000000001101";	-- 0x0AC4
		when 001379 => D <= "0110011100000000";	-- 0x0AC6
		when 001380 => D <= "0000000001100010";	-- 0x0AC8
		when 001381 => D <= "1011000111111100";	-- 0x0ACA
		when 001382 => D <= "0000000000000001";	-- 0x0ACC
		when 001383 => D <= "0000000001111111";	-- 0x0ACE
		when 001384 => D <= "0110010111000110";	-- 0x0AD0
		when 001385 => D <= "0001000000111100";	-- 0x0AD2
		when 001386 => D <= "0000000000001000";	-- 0x0AD4
		when 001387 => D <= "0110000100000000";	-- 0x0AD6
		when 001388 => D <= "1111011000110100";	-- 0x0AD8
		when 001389 => D <= "0001000000111100";	-- 0x0ADA
		when 001390 => D <= "0000000000100000";	-- 0x0ADC
		when 001391 => D <= "0110000100000000";	-- 0x0ADE
		when 001392 => D <= "1111011000101100";	-- 0x0AE0
		when 001393 => D <= "1011000111111100";	-- 0x0AE2
		when 001394 => D <= "0000000000000001";	-- 0x0AE4
		when 001395 => D <= "0000000000110000";	-- 0x0AE6
		when 001396 => D <= "0110001110101110";	-- 0x0AE8
		when 001397 => D <= "0001000000111100";	-- 0x0AEA
		when 001398 => D <= "0000000000001000";	-- 0x0AEC
		when 001399 => D <= "0110000100000000";	-- 0x0AEE
		when 001400 => D <= "1111011000011100";	-- 0x0AF0
		when 001401 => D <= "0101001110001000";	-- 0x0AF2
		when 001402 => D <= "0110000010100010";	-- 0x0AF4
		when 001403 => D <= "0010001000001000";	-- 0x0AF6
		when 001404 => D <= "0000010010000001";	-- 0x0AF8
		when 001405 => D <= "0000000000000001";	-- 0x0AFA
		when 001406 => D <= "0000000000110000";	-- 0x0AFC
		when 001407 => D <= "0110011100000000";	-- 0x0AFE
		when 001408 => D <= "0000000000100000";	-- 0x0B00
		when 001409 => D <= "0101001101000001";	-- 0x0B02
		when 001410 => D <= "0001000000111100";	-- 0x0B04
		when 001411 => D <= "0000000000001000";	-- 0x0B06
		when 001412 => D <= "0110000100000000";	-- 0x0B08
		when 001413 => D <= "1111011000000010";	-- 0x0B0A
		when 001414 => D <= "0001000000111100";	-- 0x0B0C
		when 001415 => D <= "0000000000100000";	-- 0x0B0E
		when 001416 => D <= "0110000100000000";	-- 0x0B10
		when 001417 => D <= "1111010111111010";	-- 0x0B12
		when 001418 => D <= "0001000000111100";	-- 0x0B14
		when 001419 => D <= "0000000000001000";	-- 0x0B16
		when 001420 => D <= "0110000100000000";	-- 0x0B18
		when 001421 => D <= "1111010111110010";	-- 0x0B1A
		when 001422 => D <= "0101000111001001";	-- 0x0B1C
		when 001423 => D <= "1111111111100110";	-- 0x0B1E
		when 001424 => D <= "0100000111111001";	-- 0x0B20
		when 001425 => D <= "0000000000000001";	-- 0x0B22
		when 001426 => D <= "0000000000110000";	-- 0x0B24
		when 001427 => D <= "0110000000000000";	-- 0x0B26
		when 001428 => D <= "1111111101110000";	-- 0x0B28
		when 001429 => D <= "0001000000111100";	-- 0x0B2A
		when 001430 => D <= "0000000000001010";	-- 0x0B2C
		when 001431 => D <= "0110000100000000";	-- 0x0B2E
		when 001432 => D <= "1111010111011100";	-- 0x0B30
		when 001433 => D <= "0100111001110101";	-- 0x0B32
		when 001434 => D <= "1011001010111100";	-- 0x0B34
		when 001435 => D <= "0000000000000000";	-- 0x0B36
		when 001436 => D <= "1111111111111111";	-- 0x0B38
		when 001437 => D <= "0110010000000000";	-- 0x0B3A
		when 001438 => D <= "1111111101000000";	-- 0x0B3C
		when 001439 => D <= "0010001001111000";	-- 0x0B3E
		when 001440 => D <= "0000000100000000";	-- 0x0B40
		when 001441 => D <= "0010010001111001";	-- 0x0B42
		when 001442 => D <= "0000000000000001";	-- 0x0B44
		when 001443 => D <= "0000000000100100";	-- 0x0B46
		when 001444 => D <= "0101001110001010";	-- 0x0B48
		when 001445 => D <= "1011010111001001";	-- 0x0B4A
		when 001446 => D <= "0110010100000000";	-- 0x0B4C
		when 001447 => D <= "0000000000010000";	-- 0x0B4E
		when 001448 => D <= "0001010000011001";	-- 0x0B50
		when 001449 => D <= "1110000101001010";	-- 0x0B52
		when 001450 => D <= "0001010000010001";	-- 0x0B54
		when 001451 => D <= "0101001110001001";	-- 0x0B56
		when 001452 => D <= "1011010001000001";	-- 0x0B58
		when 001453 => D <= "0110010100000000";	-- 0x0B5A
		when 001454 => D <= "0000000000000100";	-- 0x0B5C
		when 001455 => D <= "0100111001110101";	-- 0x0B5E
		when 001456 => D <= "0101010010001001";	-- 0x0B60
		when 001457 => D <= "0000110000011001";	-- 0x0B62
		when 001458 => D <= "0000000000001101";	-- 0x0B64
		when 001459 => D <= "0110011011111010";	-- 0x0B66
		when 001460 => D <= "0110000011011000";	-- 0x0B68
		when 001461 => D <= "1011011111001001";	-- 0x0B6A
		when 001462 => D <= "0110011100000000";	-- 0x0B6C
		when 001463 => D <= "0000000000000110";	-- 0x0B6E
		when 001464 => D <= "0001010011011001";	-- 0x0B70
		when 001465 => D <= "0110000011110110";	-- 0x0B72
		when 001466 => D <= "0100111001110101";	-- 0x0B74
		when 001467 => D <= "1011010111001001";	-- 0x0B76
		when 001468 => D <= "0110011111111010";	-- 0x0B78
		when 001469 => D <= "0001011100100001";	-- 0x0B7A
		when 001470 => D <= "0110000011111000";	-- 0x0B7C
		when 001471 => D <= "0010110001011111";	-- 0x0B7E
		when 001472 => D <= "0010001111011111";	-- 0x0B80
		when 001473 => D <= "0000000000000001";	-- 0x0B82
		when 001474 => D <= "0000000000010000";	-- 0x0B84
		when 001475 => D <= "0110011100000000";	-- 0x0B86
		when 001476 => D <= "0000000000011010";	-- 0x0B88
		when 001477 => D <= "0010001111011111";	-- 0x0B8A
		when 001478 => D <= "0000000000000001";	-- 0x0B8C
		when 001479 => D <= "0000000000010100";	-- 0x0B8E
		when 001480 => D <= "0010001111011111";	-- 0x0B90
		when 001481 => D <= "0000000000000001";	-- 0x0B92
		when 001482 => D <= "0000000000011000";	-- 0x0B94
		when 001483 => D <= "0010001111011111";	-- 0x0B96
		when 001484 => D <= "0000000000000001";	-- 0x0B98
		when 001485 => D <= "0000000000011100";	-- 0x0B9A
		when 001486 => D <= "0010001111011111";	-- 0x0B9C
		when 001487 => D <= "0000000000000001";	-- 0x0B9E
		when 001488 => D <= "0000000000100000";	-- 0x0BA0
		when 001489 => D <= "0100111011010110";	-- 0x0BA2
		when 001490 => D <= "0010001000111001";	-- 0x0BA4
		when 001491 => D <= "0000000000000001";	-- 0x0BA6
		when 001492 => D <= "0000000000101100";	-- 0x0BA8
		when 001493 => D <= "1001001010001111";	-- 0x0BAA
		when 001494 => D <= "0110010000000000";	-- 0x0BAC
		when 001495 => D <= "1111111011000100";	-- 0x0BAE
		when 001496 => D <= "0010110001011111";	-- 0x0BB0
		when 001497 => D <= "0010001000111001";	-- 0x0BB2
		when 001498 => D <= "0000000000000001";	-- 0x0BB4
		when 001499 => D <= "0000000000010000";	-- 0x0BB6
		when 001500 => D <= "0110011100000000";	-- 0x0BB8
		when 001501 => D <= "0000000000011010";	-- 0x0BBA
		when 001502 => D <= "0010111100111001";	-- 0x0BBC
		when 001503 => D <= "0000000000000001";	-- 0x0BBE
		when 001504 => D <= "0000000000100000";	-- 0x0BC0
		when 001505 => D <= "0010111100111001";	-- 0x0BC2
		when 001506 => D <= "0000000000000001";	-- 0x0BC4
		when 001507 => D <= "0000000000011100";	-- 0x0BC6
		when 001508 => D <= "0010111100111001";	-- 0x0BC8
		when 001509 => D <= "0000000000000001";	-- 0x0BCA
		when 001510 => D <= "0000000000011000";	-- 0x0BCC
		when 001511 => D <= "0010111100111001";	-- 0x0BCE
		when 001512 => D <= "0000000000000001";	-- 0x0BD0
		when 001513 => D <= "0000000000010100";	-- 0x0BD2
		when 001514 => D <= "0010111100000001";	-- 0x0BD4
		when 001515 => D <= "0100111011010110";	-- 0x0BD6
		when 001516 => D <= "0001001000000000";	-- 0x0BD8
		when 001517 => D <= "0001000000011001";	-- 0x0BDA
		when 001518 => D <= "1011001000000000";	-- 0x0BDC
		when 001519 => D <= "0110011100000000";	-- 0x0BDE
		when 001520 => D <= "0000000000010100";	-- 0x0BE0
		when 001521 => D <= "0110000100000000";	-- 0x0BE2
		when 001522 => D <= "1111010100101000";	-- 0x0BE4
		when 001523 => D <= "1011000000111100";	-- 0x0BE6
		when 001524 => D <= "0000000000001101";	-- 0x0BE8
		when 001525 => D <= "0110011011101110";	-- 0x0BEA
		when 001526 => D <= "0001000000111100";	-- 0x0BEC
		when 001527 => D <= "0000000000001010";	-- 0x0BEE
		when 001528 => D <= "0110000100000000";	-- 0x0BF0
		when 001529 => D <= "1111010100011010";	-- 0x0BF2
		when 001530 => D <= "0100111001110101";	-- 0x0BF4
		when 001531 => D <= "0110000100000000";	-- 0x0BF6
		when 001532 => D <= "0000000011011000";	-- 0x0BF8
		when 001533 => D <= "0010001000011001";	-- 0x0BFA
		when 001534 => D <= "0001000000111100";	-- 0x0BFC
		when 001535 => D <= "0000000000100010";	-- 0x0BFE
		when 001536 => D <= "0010001001001000";	-- 0x0C00
		when 001537 => D <= "0110000111010100";	-- 0x0C02
		when 001538 => D <= "0010000001001001";	-- 0x0C04
		when 001539 => D <= "0010001001011111";	-- 0x0C06
		when 001540 => D <= "1011000000111100";	-- 0x0C08
		when 001541 => D <= "0000000000001010";	-- 0x0C0A
		when 001542 => D <= "0110011100000000";	-- 0x0C0C
		when 001543 => D <= "1111011101101110";	-- 0x0C0E
		when 001544 => D <= "0101010010001001";	-- 0x0C10
		when 001545 => D <= "0100111011010001";	-- 0x0C12
		when 001546 => D <= "0110000100000000";	-- 0x0C14
		when 001547 => D <= "0000000010111010";	-- 0x0C16
		when 001548 => D <= "0010011100000111";	-- 0x0C18
		when 001549 => D <= "0001000000111100";	-- 0x0C1A
		when 001550 => D <= "0000000000100111";	-- 0x0C1C
		when 001551 => D <= "0110000011100000";	-- 0x0C1E
		when 001552 => D <= "0110000100000000";	-- 0x0C20
		when 001553 => D <= "0000000010101110";	-- 0x0C22
		when 001554 => D <= "0101111100001101";	-- 0x0C24
		when 001555 => D <= "0001000000111100";	-- 0x0C26
		when 001556 => D <= "0000000000001101";	-- 0x0C28
		when 001557 => D <= "0110000100000000";	-- 0x0C2A
		when 001558 => D <= "1111010011100000";	-- 0x0C2C
		when 001559 => D <= "0010001001011111";	-- 0x0C2E
		when 001560 => D <= "0110000011011110";	-- 0x0C30
		when 001561 => D <= "0100111001110101";	-- 0x0C32
		when 001562 => D <= "0010011000000001";	-- 0x0C34
		when 001563 => D <= "0011111100000100";	-- 0x0C36
		when 001564 => D <= "0001111100111100";	-- 0x0C38
		when 001565 => D <= "0000000011111111";	-- 0x0C3A
		when 001566 => D <= "0100101010000001";	-- 0x0C3C
		when 001567 => D <= "0110101000000000";	-- 0x0C3E
		when 001568 => D <= "0000000000000110";	-- 0x0C40
		when 001569 => D <= "0100010010000001";	-- 0x0C42
		when 001570 => D <= "0101001101000100";	-- 0x0C44
		when 001571 => D <= "1000001011111100";	-- 0x0C46
		when 001572 => D <= "0000000000001010";	-- 0x0C48
		when 001573 => D <= "0110100100000000";	-- 0x0C4A
		when 001574 => D <= "0000000000001110";	-- 0x0C4C
		when 001575 => D <= "0010000000000001";	-- 0x0C4E
		when 001576 => D <= "1100001010111100";	-- 0x0C50
		when 001577 => D <= "0000000000000000";	-- 0x0C52
		when 001578 => D <= "1111111111111111";	-- 0x0C54
		when 001579 => D <= "0110000000000000";	-- 0x0C56
		when 001580 => D <= "0000000000011100";	-- 0x0C58
		when 001581 => D <= "0011000000000001";	-- 0x0C5A
		when 001582 => D <= "0100001001000001";	-- 0x0C5C
		when 001583 => D <= "0100100001000001";	-- 0x0C5E
		when 001584 => D <= "1000001011111100";	-- 0x0C60
		when 001585 => D <= "0000000000001010";	-- 0x0C62
		when 001586 => D <= "0011010000000001";	-- 0x0C64
		when 001587 => D <= "0011001000000000";	-- 0x0C66
		when 001588 => D <= "1000001011111100";	-- 0x0C68
		when 001589 => D <= "0000000000001010";	-- 0x0C6A
		when 001590 => D <= "0010000000000001";	-- 0x0C6C
		when 001591 => D <= "0100100001000001";	-- 0x0C6E
		when 001592 => D <= "0011001000000010";	-- 0x0C70
		when 001593 => D <= "0100100001000001";	-- 0x0C72
		when 001594 => D <= "0100100001000000";	-- 0x0C74
		when 001595 => D <= "0001111100000000";	-- 0x0C76
		when 001596 => D <= "0100100001000000";	-- 0x0C78
		when 001597 => D <= "0101001101000100";	-- 0x0C7A
		when 001598 => D <= "0100101010000001";	-- 0x0C7C
		when 001599 => D <= "0110011011000110";	-- 0x0C7E
		when 001600 => D <= "0101001101000100";	-- 0x0C80
		when 001601 => D <= "0110101100000000";	-- 0x0C82
		when 001602 => D <= "0000000000001110";	-- 0x0C84
		when 001603 => D <= "0001000000111100";	-- 0x0C86
		when 001604 => D <= "0000000000100000";	-- 0x0C88
		when 001605 => D <= "0110000100000000";	-- 0x0C8A
		when 001606 => D <= "1111010010000000";	-- 0x0C8C
		when 001607 => D <= "0101000111001100";	-- 0x0C8E
		when 001608 => D <= "1111111111110110";	-- 0x0C90
		when 001609 => D <= "0100101010000011";	-- 0x0C92
		when 001610 => D <= "0110101000000000";	-- 0x0C94
		when 001611 => D <= "0000000000001010";	-- 0x0C96
		when 001612 => D <= "0001000000111100";	-- 0x0C98
		when 001613 => D <= "0000000000101101";	-- 0x0C9A
		when 001614 => D <= "0110000100000000";	-- 0x0C9C
		when 001615 => D <= "1111010001101110";	-- 0x0C9E
		when 001616 => D <= "0001000000011111";	-- 0x0CA0
		when 001617 => D <= "0110101100000000";	-- 0x0CA2
		when 001618 => D <= "0000000000001100";	-- 0x0CA4
		when 001619 => D <= "0000011000000000";	-- 0x0CA6
		when 001620 => D <= "0000000000110000";	-- 0x0CA8
		when 001621 => D <= "0110000100000000";	-- 0x0CAA
		when 001622 => D <= "1111010001100000";	-- 0x0CAC
		when 001623 => D <= "0110000011110000";	-- 0x0CAE
		when 001624 => D <= "0011100000011111";	-- 0x0CB0
		when 001625 => D <= "0100111001110101";	-- 0x0CB2
		when 001626 => D <= "0100001010000001";	-- 0x0CB4
		when 001627 => D <= "0001001000011001";	-- 0x0CB6
		when 001628 => D <= "1110000101001001";	-- 0x0CB8
		when 001629 => D <= "0001001000011001";	-- 0x0CBA
		when 001630 => D <= "0111100000000101";	-- 0x0CBC
		when 001631 => D <= "0110000100000000";	-- 0x0CBE
		when 001632 => D <= "1111111101110100";	-- 0x0CC0
		when 001633 => D <= "0001000000111100";	-- 0x0CC2
		when 001634 => D <= "0000000000100000";	-- 0x0CC4
		when 001635 => D <= "0110000100000000";	-- 0x0CC6
		when 001636 => D <= "1111010001000100";	-- 0x0CC8
		when 001637 => D <= "0100001001000000";	-- 0x0CCA
		when 001638 => D <= "0110000000000000";	-- 0x0CCC
		when 001639 => D <= "1111111100001010";	-- 0x0CCE
		when 001640 => D <= "0110000100000000";	-- 0x0CD0
		when 001641 => D <= "0000000001010110";	-- 0x0CD2
		when 001642 => D <= "0010001001011111";	-- 0x0CD4
		when 001643 => D <= "0001001000011001";	-- 0x0CD6
		when 001644 => D <= "1011001000010000";	-- 0x0CD8
		when 001645 => D <= "0110011100000000";	-- 0x0CDA
		when 001646 => D <= "0000000000001010";	-- 0x0CDC
		when 001647 => D <= "0100001010000001";	-- 0x0CDE
		when 001648 => D <= "0001001000010001";	-- 0x0CE0
		when 001649 => D <= "1101001111000001";	-- 0x0CE2
		when 001650 => D <= "0100111011010001";	-- 0x0CE4
		when 001651 => D <= "0101001010001000";	-- 0x0CE6
		when 001652 => D <= "0101001010001001";	-- 0x0CE8
		when 001653 => D <= "0100111011010001";	-- 0x0CEA
		when 001654 => D <= "0100001010000001";	-- 0x0CEC
		when 001655 => D <= "0100001001000010";	-- 0x0CEE
		when 001656 => D <= "0110000100000000";	-- 0x0CF0
		when 001657 => D <= "0000000000110110";	-- 0x0CF2
		when 001658 => D <= "0000110000010000";	-- 0x0CF4
		when 001659 => D <= "0000000000110000";	-- 0x0CF6
		when 001660 => D <= "0110010100000000";	-- 0x0CF8
		when 001661 => D <= "0000000000101100";	-- 0x0CFA
		when 001662 => D <= "0000110000010000";	-- 0x0CFC
		when 001663 => D <= "0000000000111001";	-- 0x0CFE
		when 001664 => D <= "0110001000000000";	-- 0x0D00
		when 001665 => D <= "0000000000100100";	-- 0x0D02
		when 001666 => D <= "1011001010111100";	-- 0x0D04
		when 001667 => D <= "0000110011001100";	-- 0x0D06
		when 001668 => D <= "1100110011001100";	-- 0x0D08
		when 001669 => D <= "0110010000000000";	-- 0x0D0A
		when 001670 => D <= "1111110101110000";	-- 0x0D0C
		when 001671 => D <= "0010000000000001";	-- 0x0D0E
		when 001672 => D <= "1101001010000001";	-- 0x0D10
		when 001673 => D <= "1101001010000001";	-- 0x0D12
		when 001674 => D <= "1101001010000000";	-- 0x0D14
		when 001675 => D <= "1101001010000001";	-- 0x0D16
		when 001676 => D <= "0001000000011000";	-- 0x0D18
		when 001677 => D <= "1100000010111100";	-- 0x0D1A
		when 001678 => D <= "0000000000000000";	-- 0x0D1C
		when 001679 => D <= "0000000000001111";	-- 0x0D1E
		when 001680 => D <= "1101001010000000";	-- 0x0D20
		when 001681 => D <= "0101001001000010";	-- 0x0D22
		when 001682 => D <= "0110000011001110";	-- 0x0D24
		when 001683 => D <= "0100111001110101";	-- 0x0D26
		when 001684 => D <= "0000110000010000";	-- 0x0D28
		when 001685 => D <= "0000000000100000";	-- 0x0D2A
		when 001686 => D <= "0110011000000000";	-- 0x0D2C
		when 001687 => D <= "0000000000000110";	-- 0x0D2E
		when 001688 => D <= "0101001010001000";	-- 0x0D30
		when 001689 => D <= "0110000011110100";	-- 0x0D32
		when 001690 => D <= "0100111001110101";	-- 0x0D34
		when 001691 => D <= "0100000111111001";	-- 0x0D36
		when 001692 => D <= "0000000000000001";	-- 0x0D38
		when 001693 => D <= "0000000000110000";	-- 0x0D3A
		when 001694 => D <= "0100001000000001";	-- 0x0D3C
		when 001695 => D <= "0001000000011000";	-- 0x0D3E
		when 001696 => D <= "1011000000111100";	-- 0x0D40
		when 001697 => D <= "0000000000001101";	-- 0x0D42
		when 001698 => D <= "0110011100000000";	-- 0x0D44
		when 001699 => D <= "0000000000100000";	-- 0x0D46
		when 001700 => D <= "1011000000111100";	-- 0x0D48
		when 001701 => D <= "0000000000100010";	-- 0x0D4A
		when 001702 => D <= "0110011100000000";	-- 0x0D4C
		when 001703 => D <= "0000000000011010";	-- 0x0D4E
		when 001704 => D <= "1011000000111100";	-- 0x0D50
		when 001705 => D <= "0000000000100111";	-- 0x0D52
		when 001706 => D <= "0110011100000000";	-- 0x0D54
		when 001707 => D <= "0000000000010010";	-- 0x0D56
		when 001708 => D <= "0100101000000001";	-- 0x0D58
		when 001709 => D <= "0110011011100010";	-- 0x0D5A
		when 001710 => D <= "0110000100000000";	-- 0x0D5C
		when 001711 => D <= "0000000000011100";	-- 0x0D5E
		when 001712 => D <= "0001000100000000";	-- 0x0D60
		when 001713 => D <= "0101001010001000";	-- 0x0D62
		when 001714 => D <= "0110000011011000";	-- 0x0D64
		when 001715 => D <= "0100111001110101";	-- 0x0D66
		when 001716 => D <= "0100101000000001";	-- 0x0D68
		when 001717 => D <= "0110011000000000";	-- 0x0D6A
		when 001718 => D <= "0000000000000110";	-- 0x0D6C
		when 001719 => D <= "0001001000000000";	-- 0x0D6E
		when 001720 => D <= "0110000011001100";	-- 0x0D70
		when 001721 => D <= "1011001000000000";	-- 0x0D72
		when 001722 => D <= "0110011011001000";	-- 0x0D74
		when 001723 => D <= "0100001000000001";	-- 0x0D76
		when 001724 => D <= "0110000011000100";	-- 0x0D78
		when 001725 => D <= "1011000000111100";	-- 0x0D7A
		when 001726 => D <= "0000000001100001";	-- 0x0D7C
		when 001727 => D <= "0110010100000000";	-- 0x0D7E
		when 001728 => D <= "0000000000001110";	-- 0x0D80
		when 001729 => D <= "1011000000111100";	-- 0x0D82
		when 001730 => D <= "0000000001111010";	-- 0x0D84
		when 001731 => D <= "0110001000000000";	-- 0x0D86
		when 001732 => D <= "0000000000000110";	-- 0x0D88
		when 001733 => D <= "0000010000000000";	-- 0x0D8A
		when 001734 => D <= "0000000000100000";	-- 0x0D8C
		when 001735 => D <= "0100111001110101";	-- 0x0D8E
		when 001736 => D <= "0110000100000000";	-- 0x0D90
		when 001737 => D <= "1111001101111110";	-- 0x0D92
		when 001738 => D <= "0110011100000000";	-- 0x0D94
		when 001739 => D <= "0000000000001110";	-- 0x0D96
		when 001740 => D <= "1011000000111100";	-- 0x0D98
		when 001741 => D <= "0000000000000011";	-- 0x0D9A
		when 001742 => D <= "0110011000000000";	-- 0x0D9C
		when 001743 => D <= "0000000000000110";	-- 0x0D9E
		when 001744 => D <= "0110000000000000";	-- 0x0DA0
		when 001745 => D <= "1111001110111010";	-- 0x0DA2
		when 001746 => D <= "0100111001110101";	-- 0x0DA4
		when 001747 => D <= "0100110111111001";	-- 0x0DA6
		when 001748 => D <= "0000000000000000";	-- 0x0DA8
		when 001749 => D <= "0000111001010110";	-- 0x0DAA
		when 001750 => D <= "0001000000011110";	-- 0x0DAC
		when 001751 => D <= "0110011100000000";	-- 0x0DAE
		when 001752 => D <= "0000000000001000";	-- 0x0DB0
		when 001753 => D <= "0110000100000000";	-- 0x0DB2
		when 001754 => D <= "1111001101011000";	-- 0x0DB4
		when 001755 => D <= "0110000011110100";	-- 0x0DB6
		when 001756 => D <= "0100111001110101";	-- 0x0DB8
		when 001757 => D <= "0000100000111001";	-- 0x0DBA
		when 001758 => D <= "0000000000000011";	-- 0x0DBC
		when 001759 => D <= "0000000000001000";	-- 0x0DBE
		when 001760 => D <= "0000000000000010";	-- 0x0DC0
		when 001761 => D <= "0110011111110110";	-- 0x0DC2
		when 001762 => D <= "0001001111000000";	-- 0x0DC4
		when 001763 => D <= "0000000000001000";	-- 0x0DC6
		when 001764 => D <= "0000000000000000";	-- 0x0DC8
		when 001765 => D <= "0100111001110101";	-- 0x0DCA
		when 001766 => D <= "0000100000111001";	-- 0x0DCC
		when 001767 => D <= "0000000000000000";	-- 0x0DCE
		when 001768 => D <= "0000000000001000";	-- 0x0DD0
		when 001769 => D <= "0000000000000010";	-- 0x0DD2
		when 001770 => D <= "0110011100000000";	-- 0x0DD4
		when 001771 => D <= "0000000000001100";	-- 0x0DD6
		when 001772 => D <= "0001000000111001";	-- 0x0DD8
		when 001773 => D <= "0000000000001000";	-- 0x0DDA
		when 001774 => D <= "0000000000000000";	-- 0x0DDC
		when 001775 => D <= "1100000000111100";	-- 0x0DDE
		when 001776 => D <= "0000000001111111";	-- 0x0DE0
		when 001777 => D <= "0100111001110101";	-- 0x0DE2
		when 001778 => D <= "0000100000111001";	-- 0x0DE4
		when 001779 => D <= "0000000000000001";	-- 0x0DE6
		when 001780 => D <= "0000000000000001";	-- 0x0DE8
		when 001781 => D <= "0000000001000001";	-- 0x0DEA
		when 001782 => D <= "0110011111110110";	-- 0x0DEC
		when 001783 => D <= "0001001111000000";	-- 0x0DEE
		when 001784 => D <= "0000000000000001";	-- 0x0DF0
		when 001785 => D <= "0000000001000011";	-- 0x0DF2
		when 001786 => D <= "0100111001110101";	-- 0x0DF4
		when 001787 => D <= "0000100000111001";	-- 0x0DF6
		when 001788 => D <= "0000000000000000";	-- 0x0DF8
		when 001789 => D <= "0000000000000001";	-- 0x0DFA
		when 001790 => D <= "0000000001000001";	-- 0x0DFC
		when 001791 => D <= "0110011100000000";	-- 0x0DFE
		when 001792 => D <= "0000000000001100";	-- 0x0E00
		when 001793 => D <= "0001000000111001";	-- 0x0E02
		when 001794 => D <= "0000000000000001";	-- 0x0E04
		when 001795 => D <= "0000000001000011";	-- 0x0E06
		when 001796 => D <= "1100000000111100";	-- 0x0E08
		when 001797 => D <= "0000000001111111";	-- 0x0E0A
		when 001798 => D <= "0100111001110101";	-- 0x0E0C
		when 001799 => D <= "0001111000111100";	-- 0x0E0E
		when 001800 => D <= "0000000011100100";	-- 0x0E10
		when 001801 => D <= "0100111001001110";	-- 0x0E12
		when 001802 => D <= "0000110100001010";	-- 0x0E14
		when 001803 => D <= "0100011101101111";	-- 0x0E16
		when 001804 => D <= "0111001001100100";	-- 0x0E18
		when 001805 => D <= "0110111100100111";	-- 0x0E1A
		when 001806 => D <= "0111001100100000";	-- 0x0E1C
		when 001807 => D <= "0100110101000011";	-- 0x0E1E
		when 001808 => D <= "0011011000111000";	-- 0x0E20
		when 001809 => D <= "0011000000110000";	-- 0x0E22
		when 001810 => D <= "0011000000100000";	-- 0x0E24
		when 001811 => D <= "0101010001101001";	-- 0x0E26
		when 001812 => D <= "0110111001111001";	-- 0x0E28
		when 001813 => D <= "0010000001000010";	-- 0x0E2A
		when 001814 => D <= "0100000101010011";	-- 0x0E2C
		when 001815 => D <= "0100100101000011";	-- 0x0E2E
		when 001816 => D <= "0010110000100000";	-- 0x0E30
		when 001817 => D <= "0111011000110001";	-- 0x0E32
		when 001818 => D <= "0010111000110010";	-- 0x0E34
		when 001819 => D <= "0000110100001010";	-- 0x0E36
		when 001820 => D <= "0000101000000000";	-- 0x0E38
		when 001821 => D <= "0000110100001010";	-- 0x0E3A
		when 001822 => D <= "0100111101001011";	-- 0x0E3C
		when 001823 => D <= "0000110100001010";	-- 0x0E3E
		when 001824 => D <= "0000000001001000";	-- 0x0E40
		when 001825 => D <= "0110111101110111";	-- 0x0E42
		when 001826 => D <= "0011111100001101";	-- 0x0E44
		when 001827 => D <= "0000101000000000";	-- 0x0E46
		when 001828 => D <= "0101011101101000";	-- 0x0E48
		when 001829 => D <= "0110000101110100";	-- 0x0E4A
		when 001830 => D <= "0011111100001101";	-- 0x0E4C
		when 001831 => D <= "0000101000000000";	-- 0x0E4E
		when 001832 => D <= "0101001101101111";	-- 0x0E50
		when 001833 => D <= "0111001001110010";	-- 0x0E52
		when 001834 => D <= "0111100100101110";	-- 0x0E54
		when 001835 => D <= "0000110100001010";	-- 0x0E56
		when 001836 => D <= "0000000000000000";	-- 0x0E58
		when others => D <= "----------------";
		end case;
	end process;
end;
